* NGSPICE file created from cap_bsw.ext - technology: sky130A

.subckt sky130_fd_pr__cap_mim_m3_1_VCTT89 m3_n386_n240# c1_n346_n200#
X0 c1_n346_n200# m3_n386_n240# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
.ends

.subckt cap_bsw VPBT1 VNBT1 VPBT2 VPBT3 VNBT3 CLKS
Xsky130_fd_pr__cap_mim_m3_1_VCTT89_0 VNBT3 VPBT3 sky130_fd_pr__cap_mim_m3_1_VCTT89
Xsky130_fd_pr__cap_mim_m3_1_VCTT89_1 VNBT3 VPBT3 sky130_fd_pr__cap_mim_m3_1_VCTT89
XXC1 VNBT1 VPBT1 sky130_fd_pr__cap_mim_m3_1_VCTT89
XXC2 CLKS VPBT2 sky130_fd_pr__cap_mim_m3_1_VCTT89
.ends

