magic
tech sky130A
magscale 1 2
timestamp 1730741762
<< pwell >>
rect -503 -3662 879 -2886
<< ndiff >>
rect -186 -3172 -134 -3120
rect 598 -3172 650 -3120
rect 510 -3427 562 -3375
<< psubdiff >>
rect -467 -2956 -365 -2922
rect 741 -2956 843 -2922
rect -467 -3096 -433 -2956
rect 809 -3096 843 -2956
rect -467 -3592 -433 -3452
rect 809 -3592 843 -3452
rect -467 -3626 -365 -3592
rect 741 -3626 843 -3592
<< psubdiffcont >>
rect -365 -2956 741 -2922
rect -467 -3452 -433 -3096
rect 809 -3452 843 -3096
rect -365 -3626 741 -3592
<< poly >>
rect 335 -3024 401 -3008
rect 335 -3058 351 -3024
rect 385 -3058 401 -3024
rect 335 -3074 401 -3058
rect 529 -3024 595 -3009
rect 529 -3058 545 -3024
rect 579 -3058 595 -3024
rect 529 -3075 595 -3058
rect 653 -3024 719 -3008
rect 653 -3058 669 -3024
rect 703 -3058 719 -3024
rect 653 -3074 719 -3058
rect -343 -3234 -277 -3218
rect -343 -3268 -327 -3234
rect -293 -3268 -277 -3234
rect -343 -3284 -277 -3268
rect -219 -3234 -153 -3218
rect -219 -3268 -203 -3234
rect -169 -3268 -153 -3234
rect -219 -3284 -153 -3268
rect -19 -3234 47 -3218
rect -19 -3268 -3 -3234
rect 31 -3268 47 -3234
rect -19 -3284 47 -3268
rect 99 -3234 159 -3222
rect 99 -3268 112 -3234
rect 146 -3268 159 -3234
rect 99 -3326 159 -3268
rect 217 -3280 277 -3222
rect 217 -3314 230 -3280
rect 264 -3314 277 -3280
rect 217 -3326 277 -3314
rect 329 -3280 395 -3264
rect 329 -3314 345 -3280
rect 379 -3314 395 -3280
rect 329 -3330 395 -3314
rect 529 -3280 595 -3264
rect 529 -3314 545 -3280
rect 579 -3314 595 -3280
rect 529 -3330 595 -3314
rect 653 -3280 719 -3264
rect 653 -3314 669 -3280
rect 703 -3314 719 -3280
rect 653 -3330 719 -3314
rect -343 -3490 -277 -3474
rect -343 -3524 -327 -3490
rect -293 -3524 -277 -3490
rect -343 -3540 -277 -3524
rect -219 -3490 -153 -3474
rect -219 -3524 -203 -3490
rect -169 -3524 -153 -3490
rect -219 -3540 -153 -3524
rect -25 -3490 41 -3474
rect -25 -3524 -9 -3490
rect 25 -3524 41 -3490
rect -25 -3540 41 -3524
<< polycont >>
rect 351 -3058 385 -3024
rect 545 -3058 579 -3024
rect 669 -3058 703 -3024
rect -327 -3268 -293 -3234
rect -203 -3268 -169 -3234
rect -3 -3268 31 -3234
rect 112 -3268 146 -3234
rect 230 -3314 264 -3280
rect 345 -3314 379 -3280
rect 545 -3314 579 -3280
rect 669 -3314 703 -3280
rect -327 -3524 -293 -3490
rect -203 -3524 -169 -3490
rect -9 -3524 25 -3490
<< locali >>
rect -467 -2956 -365 -2922
rect 741 -2956 843 -2922
rect -467 -3096 -433 -2956
rect 53 -3058 351 -3024
rect 385 -3058 441 -3024
rect 529 -3058 545 -3024
rect 579 -3058 595 -3024
rect 653 -3058 669 -3024
rect 703 -3058 729 -3024
rect -353 -3096 -231 -3062
rect 53 -3095 87 -3058
rect 289 -3108 323 -3058
rect 407 -3108 441 -3058
rect 695 -3095 729 -3058
rect 809 -3096 843 -2956
rect 689 -3196 809 -3096
rect -353 -3234 -319 -3199
rect 289 -3230 441 -3196
rect 607 -3230 729 -3196
rect -353 -3268 -327 -3234
rect -293 -3268 -277 -3234
rect -219 -3275 -203 -3234
rect -169 -3241 -3 -3234
rect -132 -3268 -3 -3241
rect 31 -3268 112 -3234
rect 146 -3264 255 -3234
rect 146 -3268 595 -3264
rect -132 -3272 595 -3268
rect -132 -3275 513 -3272
rect -219 -3280 513 -3275
rect -219 -3284 230 -3280
rect 121 -3314 230 -3284
rect 264 -3314 345 -3280
rect 379 -3306 513 -3280
rect 584 -3306 595 -3272
rect 379 -3314 545 -3306
rect 579 -3314 595 -3306
rect 653 -3314 669 -3280
rect 703 -3314 729 -3280
rect -353 -3352 -231 -3318
rect -65 -3352 87 -3318
rect 695 -3349 729 -3314
rect -433 -3452 -313 -3352
rect -467 -3592 -433 -3452
rect -353 -3490 -319 -3456
rect -65 -3490 -31 -3456
rect 53 -3490 87 -3456
rect 289 -3490 323 -3456
rect 607 -3486 729 -3452
rect -353 -3524 -327 -3490
rect -293 -3524 -277 -3490
rect -219 -3524 -211 -3490
rect -169 -3524 -153 -3490
rect -65 -3524 -9 -3490
rect 25 -3524 323 -3490
rect 809 -3592 843 -3452
rect -467 -3626 -365 -3592
rect 741 -3626 843 -3592
<< viali >>
rect 545 -3058 579 -3024
rect -327 -3268 -293 -3234
rect -203 -3268 -169 -3241
rect -169 -3268 -132 -3241
rect -203 -3275 -132 -3268
rect 513 -3280 584 -3272
rect 513 -3306 545 -3280
rect 545 -3306 579 -3280
rect 579 -3306 584 -3280
rect 669 -3314 703 -3280
rect -211 -3524 -203 -3490
rect -203 -3524 -177 -3490
<< metal1 >>
rect -279 -3068 -273 -3016
rect -221 -3030 -215 -3016
rect 539 -3024 585 -3018
rect 533 -3030 545 -3024
rect -221 -3058 545 -3030
rect 579 -3058 591 -3024
rect -221 -3068 -215 -3058
rect 539 -3064 585 -3058
rect -183 -3114 -25 -3096
rect -186 -3118 -25 -3114
rect -186 -3170 -130 -3118
rect -78 -3170 -25 -3118
rect -186 -3178 -25 -3170
rect 44 -3120 96 -3114
rect 44 -3178 96 -3172
rect 162 -3120 214 -3114
rect 162 -3178 214 -3172
rect 280 -3120 332 -3114
rect 280 -3178 332 -3172
rect 506 -3120 562 -3114
rect 558 -3172 562 -3120
rect 506 -3178 562 -3172
rect -183 -3196 -25 -3178
rect -359 -3234 -287 -3228
rect -359 -3268 -327 -3234
rect -293 -3268 -281 -3234
rect -209 -3241 -126 -3229
rect -359 -3274 -287 -3268
rect -359 -3280 -295 -3274
rect -209 -3275 -203 -3241
rect -132 -3275 -126 -3241
rect -209 -3287 -126 -3275
rect 507 -3272 590 -3260
rect 507 -3306 513 -3272
rect 584 -3306 590 -3272
rect 507 -3318 590 -3306
rect 651 -3280 715 -3262
rect 651 -3314 669 -3280
rect 703 -3314 715 -3280
rect 663 -3320 709 -3314
rect -182 -3378 -130 -3372
rect -182 -3436 -130 -3430
rect 44 -3375 96 -3369
rect 44 -3433 96 -3427
rect 162 -3375 214 -3369
rect 162 -3433 214 -3427
rect 280 -3375 283 -3369
rect 311 -3375 332 -3369
rect 280 -3433 332 -3427
rect 401 -3375 559 -3352
rect 401 -3427 454 -3375
rect 506 -3427 559 -3375
rect 401 -3452 559 -3427
rect 401 -3480 429 -3452
rect -279 -3532 -273 -3480
rect -221 -3490 -165 -3480
rect -221 -3524 -211 -3490
rect -177 -3524 -165 -3490
rect -221 -3532 -165 -3524
rect -136 -3532 -130 -3480
rect -78 -3508 429 -3480
rect -78 -3532 -72 -3508
<< via1 >>
rect -273 -3068 -221 -3016
rect -130 -3170 -78 -3118
rect 44 -3172 96 -3120
rect 162 -3172 214 -3120
rect 280 -3172 332 -3120
rect 506 -3172 558 -3120
rect -182 -3430 -130 -3378
rect 44 -3427 96 -3375
rect 162 -3427 214 -3375
rect 280 -3427 332 -3375
rect 454 -3427 506 -3375
rect -273 -3532 -221 -3480
rect -130 -3532 -78 -3480
<< metal2 >>
rect -273 -3016 -221 -3010
rect -273 -3480 -221 -3068
rect -130 -3118 -78 -3112
rect -130 -3372 -78 -3170
rect -182 -3378 -78 -3372
rect -130 -3430 -78 -3378
rect -182 -3436 -78 -3430
rect 44 -3120 96 -3114
rect 44 -3375 96 -3172
rect 44 -3433 96 -3427
rect 162 -3120 214 -3114
rect 162 -3375 214 -3172
rect 162 -3433 214 -3427
rect 280 -3120 332 -3114
rect 280 -3375 332 -3172
rect 280 -3433 332 -3427
rect 454 -3375 506 -3120
rect 558 -3172 564 -3120
rect 454 -3433 506 -3427
rect -273 -3538 -221 -3532
rect -130 -3480 -78 -3436
rect -130 -3538 -78 -3532
use sky130_fd_pr__nfet_01v8_6J3TAM  sky130_fd_pr__nfet_01v8_6J3TAM_0
timestamp 1730727801
transform 1 0 -204 0 1 -3146
box -73 -76 73 76
use sky130_fd_pr__nfet_01v8_6J3TAM  sky130_fd_pr__nfet_01v8_6J3TAM_1
timestamp 1730727801
transform 1 0 580 0 1 -3402
box -73 -76 73 76
use sky130_fd_pr__nfet_01v8_6J3TAM  sky130_fd_pr__nfet_01v8_6J3TAM_2
timestamp 1730727801
transform 1 0 -204 0 1 -3402
box -73 -76 73 76
use sky130_fd_pr__nfet_01v8_6J3TAM  sky130_fd_pr__nfet_01v8_6J3TAM_3
timestamp 1730727801
transform 1 0 580 0 1 -3146
box -73 -76 73 76
use sky130_fd_pr__nfet_01v8_6J3TAM  sky130_fd_pr__nfet_01v8_6J3TAM_4
timestamp 1730727801
transform 1 0 668 0 1 -3146
box -73 -76 73 76
use sky130_fd_pr__nfet_01v8_6J3TAM  sky130_fd_pr__nfet_01v8_6J3TAM_5
timestamp 1730727801
transform 1 0 -292 0 1 -3402
box -73 -76 73 76
use sky130_fd_pr__nfet_01v8_6J3TAM  sky130_fd_pr__nfet_01v8_6J3TAM_6
timestamp 1730727801
transform 1 0 668 0 1 -3402
box -73 -76 73 76
use sky130_fd_pr__nfet_01v8_6J3TAM  sky130_fd_pr__nfet_01v8_6J3TAM_10
timestamp 1730727801
transform 1 0 -292 0 1 -3146
box -73 -76 73 76
use sky130_fd_pr__nfet_01v8_QS6TK8  sky130_fd_pr__nfet_01v8_QS6TK8_0
timestamp 1730727801
transform 1 0 11 0 1 -3146
box -88 -76 88 76
use sky130_fd_pr__nfet_01v8_QS6TK8  sky130_fd_pr__nfet_01v8_QS6TK8_1
timestamp 1730727801
transform 1 0 129 0 1 -3146
box -88 -76 88 76
use sky130_fd_pr__nfet_01v8_QS6TK8  sky130_fd_pr__nfet_01v8_QS6TK8_2
timestamp 1730727801
transform 1 0 247 0 1 -3146
box -88 -76 88 76
use sky130_fd_pr__nfet_01v8_QS6TK8  sky130_fd_pr__nfet_01v8_QS6TK8_3
timestamp 1730727801
transform 1 0 365 0 1 -3402
box -88 -76 88 76
use sky130_fd_pr__nfet_01v8_QS6TK8  sky130_fd_pr__nfet_01v8_QS6TK8_4
timestamp 1730727801
transform 1 0 365 0 1 -3146
box -88 -76 88 76
use sky130_fd_pr__nfet_01v8_QS6TK8  sky130_fd_pr__nfet_01v8_QS6TK8_5
timestamp 1730727801
transform 1 0 11 0 1 -3402
box -88 -76 88 76
use sky130_fd_pr__nfet_01v8_QS6TK8  sky130_fd_pr__nfet_01v8_QS6TK8_6
timestamp 1730727801
transform 1 0 129 0 1 -3402
box -88 -76 88 76
use sky130_fd_pr__nfet_01v8_QS6TK8  sky130_fd_pr__nfet_01v8_QS6TK8_7
timestamp 1730727801
transform 1 0 247 0 1 -3402
box -88 -76 88 76
<< labels >>
flabel metal2 s 71 -3290 71 -3290 0 FreeSans 320 0 0 0 VI
port 1 nsew
flabel metal1 s -188 -3255 -188 -3255 0 FreeSans 320 0 0 0 VBOOT
port 2 nsew
flabel metal2 s -104 -3331 -104 -3331 0 FreeSans 320 0 0 0 VNBT3
port 4 nsew
flabel metal1 s -342 -3252 -342 -3252 0 FreeSans 320 0 0 0 SWITCHING
port 5 nsew
flabel metal1 s 684 -3298 684 -3298 0 FreeSans 320 0 0 0 SWITCHING
flabel locali s 184 -2937 184 -2937 0 FreeSans 320 0 0 0 VSSA
port 6 nsew
flabel metal1 s -115 -3042 -115 -3042 0 FreeSans 320 0 0 0 VNBT1
port 3 nsew
flabel metal2 s 187 -3329 187 -3329 0 FreeSans 320 0 0 0 VO
port 7 nsew
<< end >>
