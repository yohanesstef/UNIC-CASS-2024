* NGSPICE file created from sample-n-hold-layout.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_LCNWMQ a_15_n90# a_n33_n187# w_n211_n310# a_n73_n90#
+ VSUBS
X0 a_15_n90# a_n33_n187# a_n73_n90# w_n211_n310# sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
C0 a_n73_n90# a_15_n90# 0.203436f
C1 w_n211_n310# a_n73_n90# 0.101688f
C2 a_n33_n187# a_n73_n90# 0.015928f
C3 w_n211_n310# a_15_n90# 0.101688f
C4 a_n33_n187# a_15_n90# 0.015928f
C5 w_n211_n310# a_n33_n187# 0.14302f
C6 a_15_n90# VSUBS 0.062251f
C7 a_n73_n90# VSUBS 0.062251f
C8 a_n33_n187# VSUBS 0.080068f
C9 w_n211_n310# VSUBS 1.19627f
.ends

.subckt sky130_fd_pr__nfet_01v8_L78EGD a_n33_33# a_15_n73# a_n73_n73# a_n175_n185#
X0 a_15_n73# a_n33_33# a_n73_n73# a_n175_n185# sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
C0 a_n73_n73# a_n33_33# 0.012054f
C1 a_15_n73# a_n73_n73# 0.069931f
C2 a_15_n73# a_n33_33# 0.012054f
C3 a_15_n73# a_n175_n185# 0.078869f
C4 a_n73_n73# a_n175_n185# 0.078869f
C5 a_n33_33# a_n175_n185# 0.220946f
.ends

.subckt sky130_fd_pr__nfet_01v8_TK2CNP a_30_n531# a_n33_491# a_n88_n531# a_n190_n643#
X0 a_30_n531# a_n33_491# a_n88_n531# a_n190_n643# sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=0.3
C0 a_n88_n531# a_30_n531# 0.595979f
C1 a_n33_491# a_30_n531# 0.04201f
C2 a_n88_n531# a_n33_491# 0.04201f
C3 a_30_n531# a_n190_n643# 0.555909f
C4 a_n88_n531# a_n190_n643# 0.555909f
C5 a_n33_491# a_n190_n643# 0.234139f
.ends

.subckt sky130_fd_pr__pfet_01v8_M4BBJH w_n211_n384# a_n73_n164# a_n33_n261# a_15_n164#
+ VSUBS
X0 a_15_n164# a_n33_n261# a_n73_n164# w_n211_n384# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
C0 a_n33_n261# a_15_n164# 0.019421f
C1 a_n73_n164# a_15_n164# 0.321048f
C2 w_n211_n384# a_n33_n261# 0.142016f
C3 w_n211_n384# a_n73_n164# 0.146809f
C4 w_n211_n384# a_15_n164# 0.146809f
C5 a_n33_n261# a_n73_n164# 0.019421f
C6 a_15_n164# VSUBS 0.092202f
C7 a_n73_n164# VSUBS 0.092202f
C8 a_n33_n261# VSUBS 0.07969f
C9 w_n211_n384# VSUBS 1.45693f
.ends

.subckt sky130_fd_pr__nfet_01v8_7XY3PK a_15_n131# a_n175_n243# a_n33_91# a_n73_n131#
X0 a_15_n131# a_n33_91# a_n73_n131# a_n175_n243# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 a_n73_n131# a_n33_91# 0.015495f
C1 a_15_n131# a_n73_n131# 0.162113f
C2 a_15_n131# a_n33_91# 0.015495f
C3 a_15_n131# a_n175_n243# 0.13771f
C4 a_n73_n131# a_n175_n243# 0.13771f
C5 a_n33_91# a_n175_n243# 0.218066f
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_5XYVA6 m3_n893_n747# c1_n853_n707# VSUBS
X0 c1_n853_n707# m3_n893_n747# sky130_fd_pr__cap_mim_m3_1 l=7.07 w=7.07
C0 c1_n853_n707# m3_n893_n747# 4.95002f
C1 c1_n853_n707# VSUBS 0.703986f
C2 m3_n893_n747# VSUBS 2.48364f
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_5XY9G7 m3_n893_n747# c1_n853_n707# VSUBS
X0 c1_n853_n707# m3_n893_n747# sky130_fd_pr__cap_mim_m3_1 l=7.07 w=7.07
C0 m3_n893_n747# c1_n853_n707# 4.95002f
C1 c1_n853_n707# VSUBS 0.703986f
C2 m3_n893_n747# VSUBS 2.48364f
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_QEFW4K c1_n2377_n2231# m3_n2417_n2271# VSUBS
X0 c1_n2377_n2231# m3_n2417_n2271# sky130_fd_pr__cap_mim_m3_1 l=22.31 w=22.31
C0 c1_n2377_n2231# m3_n2417_n2271# 44.3143f
C1 c1_n2377_n2231# VSUBS 2.31009f
C2 m3_n2417_n2271# VSUBS 11.5049f
.ends

.subckt sample-n-hold-layout clk vdata VDD GND Vout
XXM13 m1_n220_n322# clk VDD VDD GND sky130_fd_pr__pfet_01v8_LCNWMQ
XXM15 m1_96_n322# m1_n220_n322# VDD VDD GND sky130_fd_pr__pfet_01v8_LCNWMQ
XXM16 m1_n220_n322# m1_96_n322# GND GND sky130_fd_pr__nfet_01v8_L78EGD
Xsky130_fd_pr__nfet_01v8_L78EGD_0 clk m1_n220_n322# GND GND sky130_fd_pr__nfet_01v8_L78EGD
Xsky130_fd_pr__nfet_01v8_TK2CNP_0 Vout vboot vdata GND sky130_fd_pr__nfet_01v8_TK2CNP
Xsky130_fd_pr__pfet_01v8_LCNWMQ_0 m1_412_n322# m1_96_n322# VDD VDD GND sky130_fd_pr__pfet_01v8_LCNWMQ
XXM1 c1_up VDD m1_1333_n260# GND sky130_fd_pr__nfet_01v8_L78EGD
XXM2 c3_up c3_up m1_412_n322# vboot GND sky130_fd_pr__pfet_01v8_M4BBJH
XXM3 m1_1333_n260# VDD c1_up GND sky130_fd_pr__nfet_01v8_L78EGD
XXM4 c3_up GND c1_up VDD sky130_fd_pr__nfet_01v8_7XY3PK
XXM5 m1_n220_n322# GND m1_316_n469# GND sky130_fd_pr__nfet_01v8_L78EGD
XXM7 m1_96_n322# m1_412_n322# m1_316_n469# GND sky130_fd_pr__nfet_01v8_L78EGD
XXM9 m1_n220_n322# GND m1_2597_n322# GND sky130_fd_pr__nfet_01v8_L78EGD
XXM8 VDD m1_2597_n322# vboot GND sky130_fd_pr__nfet_01v8_L78EGD
XXC1 m1_n220_n322# c1_up GND sky130_fd_pr__cap_mim_m3_1_5XYVA6
XXC2 m1_96_n322# m1_1333_n260# GND sky130_fd_pr__cap_mim_m3_1_5XY9G7
XXC3 c3_up m1_316_n469# GND sky130_fd_pr__cap_mim_m3_1_QEFW4K
XXM10 vboot m1_316_n469# m1_412_n322# GND sky130_fd_pr__nfet_01v8_L78EGD
XXM11 vdata GND vboot m1_316_n469# sky130_fd_pr__nfet_01v8_7XY3PK
C0 vboot VDD 1.601413f
C1 VDD Vout 0.065603f
C2 VDD c3_up 2.897374f
C3 c1_up VDD 1.048535f
C4 VDD m1_316_n469# 2.127093f
C5 vboot m1_412_n322# 0.677711f
C6 m1_2597_n322# VDD 0.005684f
C7 VDD m1_n220_n322# 2.160496f
C8 VDD vdata 3.16e-19
C9 m1_412_n322# c3_up 0.60504f
C10 c1_up m1_412_n322# 0.502128f
C11 VDD m1_1333_n260# 3.132697f
C12 m1_412_n322# m1_316_n469# 0.03479f
C13 vboot m1_96_n322# 0.182125f
C14 m1_412_n322# m1_n220_n322# 0.30873f
C15 m1_96_n322# c3_up 0.344904f
C16 c1_up m1_96_n322# 0.534458f
C17 m1_412_n322# m1_1333_n260# 0.096882f
C18 m1_96_n322# m1_316_n469# 0.439068f
C19 VDD clk 0.350417f
C20 m1_96_n322# m1_n220_n322# 1.322518f
C21 m1_96_n322# m1_1333_n260# 0.611439f
C22 m1_412_n322# clk 9.1e-22
C23 vboot Vout 0.090617f
C24 vboot c3_up 0.309196f
C25 c1_up vboot 3.78e-19
C26 Vout c3_up 0.038841f
C27 c1_up c3_up 0.5849f
C28 vboot m1_316_n469# 0.441249f
C29 vboot m1_2597_n322# 0.017335f
C30 vboot m1_n220_n322# 0.41364f
C31 m1_316_n469# c3_up 0.661757f
C32 c1_up m1_316_n469# 0.39875f
C33 Vout m1_n220_n322# 2.76e-19
C34 vboot vdata 0.151728f
C35 m1_2597_n322# c3_up 0.001624f
C36 Vout vdata 0.09484f
C37 m1_n220_n322# c3_up 0.584858f
C38 c1_up m1_n220_n322# 0.712525f
C39 vboot m1_1333_n260# 0.545133f
C40 vdata c3_up 0.010764f
C41 m1_2597_n322# m1_316_n469# 0.076876f
C42 m1_n220_n322# m1_316_n469# 0.29749f
C43 m1_1333_n260# c3_up 0.482581f
C44 c1_up m1_1333_n260# 0.490845f
C45 m1_2597_n322# m1_n220_n322# 0.004666f
C46 vdata m1_316_n469# 0.053263f
C47 m1_n220_n322# vdata 2.17e-19
C48 m1_1333_n260# m1_316_n469# 0.358933f
C49 m1_2597_n322# m1_1333_n260# 4.37e-19
C50 m1_1333_n260# m1_n220_n322# 0.139157f
C51 m1_412_n322# VDD 1.057846f
C52 clk m1_n220_n322# 0.708163f
C53 m1_96_n322# VDD 1.984722f
C54 m1_96_n322# m1_412_n322# 0.896762f
C55 vdata GND 1.930537f
C56 m1_2597_n322# GND 0.238383f
C57 m1_412_n322# GND 0.911725f
C58 m1_316_n469# GND 13.832773f
C59 c1_up GND 2.565598f
C60 m1_1333_n260# GND 1.197823f
C61 vboot GND 1.642715f
C62 c3_up GND 4.409274f
C63 Vout GND 1.089422f
C64 m1_96_n322# GND 2.781989f
C65 m1_n220_n322# GND 4.561662f
C66 VDD GND 11.968059f
C67 clk GND 0.776164f
.ends

