* NGSPICE file created from sample-n-hold-layout.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_LCNWMQ a_15_n90# a_n33_n187# w_n211_n310# a_n73_n90#
+ VSUBS
X0 a_15_n90# a_n33_n187# a_n73_n90# w_n211_n310# sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
C0 w_n211_n310# a_n33_n187# 0.14302f
C1 a_n73_n90# w_n211_n310# 0.101688f
C2 w_n211_n310# a_15_n90# 0.101688f
C3 a_n73_n90# a_n33_n187# 0.015928f
C4 a_n33_n187# a_15_n90# 0.015928f
C5 a_n73_n90# a_15_n90# 0.203436f
C6 a_15_n90# VSUBS 0.062251f
C7 a_n73_n90# VSUBS 0.062251f
C8 a_n33_n187# VSUBS 0.080068f
C9 w_n211_n310# VSUBS 1.19627f
.ends

.subckt sky130_fd_pr__nfet_01v8_L78EGD a_n33_33# a_15_n73# a_n73_n73# a_n175_n185#
X0 a_15_n73# a_n33_33# a_n73_n73# a_n175_n185# sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
C0 a_n73_n73# a_15_n73# 0.069931f
C1 a_n33_33# a_n73_n73# 0.012054f
C2 a_n33_33# a_15_n73# 0.012054f
C3 a_15_n73# a_n175_n185# 0.078869f
C4 a_n73_n73# a_n175_n185# 0.078869f
C5 a_n33_33# a_n175_n185# 0.220946f
.ends

.subckt sky130_fd_pr__nfet_01v8_TK2CNP a_30_n531# a_n33_491# a_n88_n531# a_n190_n643#
X0 a_30_n531# a_n33_491# a_n88_n531# a_n190_n643# sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=0.3
C0 a_n88_n531# a_n33_491# 0.04201f
C1 a_30_n531# a_n88_n531# 0.595979f
C2 a_30_n531# a_n33_491# 0.04201f
C3 a_30_n531# a_n190_n643# 0.555909f
C4 a_n88_n531# a_n190_n643# 0.555909f
C5 a_n33_491# a_n190_n643# 0.234139f
.ends

.subckt sky130_fd_pr__pfet_01v8_M4BBJH w_n211_n384# a_n73_n164# a_n33_n261# a_15_n164#
+ VSUBS
X0 a_15_n164# a_n33_n261# a_n73_n164# w_n211_n384# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
C0 a_n33_n261# w_n211_n384# 0.142016f
C1 a_n33_n261# a_n73_n164# 0.019421f
C2 w_n211_n384# a_n73_n164# 0.146809f
C3 a_15_n164# a_n33_n261# 0.019421f
C4 a_15_n164# w_n211_n384# 0.146809f
C5 a_15_n164# a_n73_n164# 0.321048f
C6 a_15_n164# VSUBS 0.092202f
C7 a_n73_n164# VSUBS 0.092202f
C8 a_n33_n261# VSUBS 0.07969f
C9 w_n211_n384# VSUBS 1.45693f
.ends

.subckt sky130_fd_pr__nfet_01v8_7XY3PK a_15_n131# a_n175_n243# a_n33_91# a_n73_n131#
X0 a_15_n131# a_n33_91# a_n73_n131# a_n175_n243# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 a_n73_n131# a_15_n131# 0.162113f
C1 a_n33_91# a_n73_n131# 0.015495f
C2 a_n33_91# a_15_n131# 0.015495f
C3 a_15_n131# a_n175_n243# 0.13771f
C4 a_n73_n131# a_n175_n243# 0.13771f
C5 a_n33_91# a_n175_n243# 0.218066f
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_5XYVA6 m3_n893_n747# c1_n853_n707# VSUBS
X0 c1_n853_n707# m3_n893_n747# sky130_fd_pr__cap_mim_m3_1 l=7.07 w=7.07
C0 c1_n853_n707# m3_n893_n747# 4.95002f
C1 c1_n853_n707# VSUBS 0.703986f
C2 m3_n893_n747# VSUBS 2.48364f
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_5XY9G7 m3_n893_n747# c1_n853_n707# VSUBS
X0 c1_n853_n707# m3_n893_n747# sky130_fd_pr__cap_mim_m3_1 l=7.07 w=7.07
C0 c1_n853_n707# m3_n893_n747# 4.95002f
C1 c1_n853_n707# VSUBS 0.703986f
C2 m3_n893_n747# VSUBS 2.48364f
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_QEFW4K c1_n2377_n2231# m3_n2417_n2271# VSUBS
X0 c1_n2377_n2231# m3_n2417_n2271# sky130_fd_pr__cap_mim_m3_1 l=22.31 w=22.31
C0 m3_n2417_n2271# c1_n2377_n2231# 44.3143f
C1 c1_n2377_n2231# VSUBS 2.31009f
C2 m3_n2417_n2271# VSUBS 11.5049f
.ends

.subckt sample-n-hold-layout clk vdata VDD GND Vout
XXM13 m1_n220_n322# clk VDD VDD GND sky130_fd_pr__pfet_01v8_LCNWMQ
XXM15 m1_96_n322# m1_n220_n322# VDD VDD GND sky130_fd_pr__pfet_01v8_LCNWMQ
XXM16 m1_n220_n322# m1_96_n322# GND GND sky130_fd_pr__nfet_01v8_L78EGD
Xsky130_fd_pr__nfet_01v8_L78EGD_0 clk m1_n220_n322# GND GND sky130_fd_pr__nfet_01v8_L78EGD
Xsky130_fd_pr__nfet_01v8_TK2CNP_0 Vout vboot vdata GND sky130_fd_pr__nfet_01v8_TK2CNP
Xsky130_fd_pr__pfet_01v8_LCNWMQ_0 m1_412_n322# m1_96_n322# VDD VDD GND sky130_fd_pr__pfet_01v8_LCNWMQ
XXM1 m1_876_n400# VDD m1_1333_n260# GND sky130_fd_pr__nfet_01v8_L78EGD
XXM2 li_891_829# li_891_829# m1_412_n322# vboot GND sky130_fd_pr__pfet_01v8_M4BBJH
XXM3 m1_1333_n260# VDD m1_876_n400# GND sky130_fd_pr__nfet_01v8_L78EGD
XXM4 li_891_829# GND m1_876_n400# VDD sky130_fd_pr__nfet_01v8_7XY3PK
XXM5 m1_n220_n322# GND m1_316_n469# GND sky130_fd_pr__nfet_01v8_L78EGD
XXM7 m1_96_n322# m1_412_n322# m1_316_n469# GND sky130_fd_pr__nfet_01v8_L78EGD
XXM9 m1_n220_n322# GND m1_2597_n322# GND sky130_fd_pr__nfet_01v8_L78EGD
XXM8 VDD m1_2597_n322# vboot GND sky130_fd_pr__nfet_01v8_L78EGD
XXC1 m1_n220_n322# m1_876_n400# GND sky130_fd_pr__cap_mim_m3_1_5XYVA6
XXC2 m1_96_n322# m1_1333_n260# GND sky130_fd_pr__cap_mim_m3_1_5XY9G7
XXC3 li_891_829# m1_316_n469# GND sky130_fd_pr__cap_mim_m3_1_QEFW4K
XXM10 vboot m1_316_n469# m1_412_n322# GND sky130_fd_pr__nfet_01v8_L78EGD
XXM11 vdata GND vboot m1_316_n469# sky130_fd_pr__nfet_01v8_7XY3PK
C0 li_891_829# m1_412_n322# 0.465194f
C1 clk VDD 0.350417f
C2 m1_96_n322# VDD 3.354356f
C3 m1_n220_n322# VDD 2.309469f
C4 clk m1_876_n400# 0.004275f
C5 li_891_829# m1_2597_n322# 0.003633f
C6 Vout li_891_829# 0.018245f
C7 m1_96_n322# m1_876_n400# 0.74927f
C8 m1_n220_n322# m1_876_n400# 1.177665f
C9 m1_1333_n260# VDD 2.795697f
C10 vdata VDD 3.16e-19
C11 m1_96_n322# clk 0.00223f
C12 m1_n220_n322# clk 0.602611f
C13 m1_1333_n260# m1_876_n400# 0.492715f
C14 m1_96_n322# m1_n220_n322# 2.654504f
C15 vboot VDD 1.619323f
C16 m1_316_n469# VDD 0.083504f
C17 m1_1333_n260# clk 1.33e-19
C18 vboot m1_876_n400# 0.117498f
C19 m1_316_n469# m1_876_n400# 0.379745f
C20 m1_412_n322# VDD 1.078815f
C21 m1_1333_n260# m1_96_n322# 0.372644f
C22 m1_1333_n260# m1_n220_n322# 0.972581f
C23 m1_96_n322# vdata 0.042761f
C24 m1_n220_n322# vdata 2.3e-19
C25 m1_876_n400# m1_412_n322# 0.202743f
C26 vboot clk 1.03e-20
C27 m1_2597_n322# VDD 0.005684f
C28 Vout VDD 0.065603f
C29 li_891_829# VDD 1.688823f
C30 m1_96_n322# vboot 0.635864f
C31 m1_n220_n322# vboot 0.878999f
C32 m1_316_n469# m1_96_n322# 0.292326f
C33 m1_316_n469# m1_n220_n322# 0.463067f
C34 clk m1_412_n322# 1.92e-19
C35 li_891_829# m1_876_n400# 0.071188f
C36 m1_96_n322# m1_412_n322# 1.426704f
C37 m1_n220_n322# m1_412_n322# 0.982966f
C38 m1_1333_n260# vboot 0.562548f
C39 m1_1333_n260# m1_316_n469# 0.035464f
C40 vboot vdata 0.151728f
C41 li_891_829# clk 0.002356f
C42 m1_316_n469# vdata 0.1334f
C43 m1_96_n322# m1_2597_n322# 0.020565f
C44 m1_n220_n322# m1_2597_n322# 0.004666f
C45 Vout m1_96_n322# 0.041538f
C46 Vout m1_n220_n322# 2.76e-19
C47 m1_96_n322# li_891_829# 0.347884f
C48 m1_n220_n322# li_891_829# 0.78406f
C49 m1_1333_n260# m1_412_n322# 0.094732f
C50 m1_316_n469# vboot 0.351288f
C51 m1_1333_n260# m1_2597_n322# 1.38e-19
C52 vboot m1_412_n322# 0.677711f
C53 m1_1333_n260# li_891_829# 0.02271f
C54 m1_316_n469# m1_412_n322# 0.048731f
C55 Vout vdata 0.09484f
C56 li_891_829# vdata 0.035611f
C57 vboot m1_2597_n322# 0.017335f
C58 Vout vboot 0.090617f
C59 li_891_829# vboot 0.035926f
C60 m1_316_n469# m1_2597_n322# 0.083365f
C61 Vout m1_316_n469# 0.02732f
C62 m1_876_n400# VDD 0.526285f
C63 m1_316_n469# li_891_829# 0.33265f
C64 vdata GND 1.930537f
C65 vboot GND 1.697857f
C66 m1_316_n469# GND 15.177321f
C67 m1_2597_n322# GND 0.238403f
C68 m1_412_n322# GND 0.971661f
C69 li_891_829# GND 3.894805f
C70 VDD GND 11.967019f
C71 m1_876_n400# GND 1.898908f
C72 m1_1333_n260# GND 1.148744f
C73 Vout GND 1.089422f
C74 clk GND 0.776164f
C75 m1_96_n322# GND 2.660355f
C76 m1_n220_n322# GND 3.057423f
.ends

