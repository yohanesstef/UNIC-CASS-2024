magic
tech sky130A
magscale 1 2
timestamp 1730554222
<< pwell >>
rect 4653 -1676 5339 -261
<< psubdiff >>
rect 4689 -332 4791 -297
rect 5201 -332 5303 -297
rect 4689 -497 4723 -332
rect 5269 -497 5303 -332
rect 4689 -1605 4723 -1419
rect 5269 -1605 5303 -1419
rect 4689 -1640 4791 -1605
rect 5201 -1640 5303 -1605
<< psubdiffcont >>
rect 4791 -332 5201 -297
rect 4689 -1419 4723 -497
rect 5269 -1419 5303 -497
rect 4791 -1640 5201 -1605
<< poly >>
rect 4813 -379 4879 -363
rect 4813 -413 4829 -379
rect 4863 -413 4879 -379
rect 4813 -429 4879 -413
rect 4989 -379 5055 -363
rect 4989 -413 5005 -379
rect 5039 -413 5055 -379
rect 4989 -429 5055 -413
rect 4849 -471 4879 -429
rect 5025 -471 5055 -429
rect 5113 -379 5179 -363
rect 5113 -413 5129 -379
rect 5163 -413 5179 -379
rect 5113 -429 5179 -413
rect 5113 -471 5143 -429
rect 4813 -681 4879 -665
rect 4813 -715 4829 -681
rect 4863 -715 4879 -681
rect 4813 -731 4879 -715
rect 4937 -731 4967 -623
rect 5113 -681 5179 -665
rect 5113 -701 5129 -681
rect 5025 -715 5129 -701
rect 5163 -715 5179 -681
rect 5025 -731 5179 -715
rect 4937 -925 4967 -883
rect 4937 -940 5055 -925
rect 4937 -974 4953 -940
rect 5039 -974 5055 -940
rect 4937 -991 5055 -974
rect 5025 -1033 5055 -991
rect 4813 -1201 4967 -1185
rect 4813 -1235 4829 -1201
rect 4863 -1215 4967 -1201
rect 4863 -1235 4879 -1215
rect 4813 -1251 4879 -1235
rect 5025 -1293 5055 -1185
rect 5113 -1201 5179 -1185
rect 5113 -1235 5129 -1201
rect 5163 -1235 5179 -1201
rect 5113 -1251 5179 -1235
rect 4849 -1487 4879 -1419
rect 4813 -1503 4879 -1487
rect 4813 -1537 4829 -1503
rect 4863 -1537 4879 -1503
rect 4813 -1553 4879 -1537
rect 4937 -1487 4967 -1419
rect 5113 -1487 5143 -1419
rect 4937 -1503 5003 -1487
rect 4937 -1537 4953 -1503
rect 4987 -1537 5003 -1503
rect 4937 -1553 5003 -1537
rect 5113 -1503 5179 -1487
rect 5113 -1537 5129 -1503
rect 5163 -1537 5179 -1503
rect 5113 -1553 5179 -1537
<< polycont >>
rect 4829 -413 4863 -379
rect 5005 -413 5039 -379
rect 5129 -413 5163 -379
rect 4829 -715 4863 -681
rect 5129 -715 5163 -681
rect 4953 -974 5039 -940
rect 4829 -1235 4863 -1201
rect 5129 -1235 5163 -1201
rect 4829 -1537 4863 -1503
rect 4953 -1537 4987 -1503
rect 5129 -1537 5163 -1503
<< locali >>
rect 4689 -332 4791 -297
rect 5201 -332 5303 -297
rect 4689 -497 4723 -332
rect 4813 -413 4829 -379
rect 4863 -413 4879 -379
rect 4989 -413 5005 -379
rect 5039 -413 5055 -379
rect 5113 -413 5129 -379
rect 5163 -413 5179 -379
rect 5269 -497 5303 -332
rect 4813 -715 4829 -681
rect 4863 -715 4879 -681
rect 5113 -715 5129 -681
rect 5163 -715 5179 -681
rect 4839 -974 4953 -940
rect 5039 -974 5154 -940
rect 4813 -1235 4829 -1201
rect 4863 -1235 4879 -1201
rect 5113 -1235 5129 -1201
rect 5163 -1235 5179 -1201
rect 4689 -1605 4723 -1419
rect 4813 -1537 4829 -1503
rect 4863 -1537 4879 -1503
rect 4937 -1537 4953 -1503
rect 4987 -1537 5003 -1503
rect 5113 -1537 5129 -1503
rect 5163 -1537 5179 -1503
rect 5269 -1605 5303 -1419
rect 4689 -1640 4791 -1605
rect 5201 -1640 5303 -1605
<< viali >>
rect 4829 -413 4863 -379
rect 5005 -413 5039 -379
rect 5129 -413 5163 -379
rect 4829 -715 4863 -681
rect 5129 -715 5163 -681
rect 4805 -974 4839 -940
rect 5154 -974 5188 -940
rect 4829 -1235 4863 -1201
rect 5129 -1235 5163 -1201
rect 4829 -1537 4863 -1503
rect 4953 -1537 4987 -1503
rect 5129 -1537 5163 -1503
<< metal1 >>
rect 4995 -371 5047 -363
rect 4815 -379 4875 -373
rect 4815 -413 4829 -379
rect 4863 -391 4875 -379
rect 4993 -377 5051 -371
rect 4993 -391 4994 -377
rect 4863 -413 4994 -391
rect 4815 -419 4994 -413
rect 4815 -509 4843 -419
rect 4903 -497 4931 -419
rect 4993 -429 4994 -419
rect 5046 -419 5051 -377
rect 5117 -379 5177 -373
rect 5117 -391 5129 -379
rect 5079 -413 5129 -391
rect 5163 -413 5177 -379
rect 5079 -419 5177 -413
rect 5046 -429 5047 -419
rect 4994 -435 5046 -429
rect 5079 -497 5107 -419
rect 5149 -497 5177 -419
rect 5058 -523 5110 -517
rect 5058 -581 5110 -575
rect 4823 -681 4869 -669
rect 4823 -699 4829 -681
rect 4815 -715 4829 -699
rect 4863 -699 4869 -681
rect 4973 -675 5019 -597
rect 4973 -681 5177 -675
rect 4863 -715 4913 -699
rect 4815 -727 4913 -715
rect 4815 -758 4843 -727
rect 4885 -757 4913 -727
rect 4973 -715 5129 -681
rect 5163 -715 5177 -681
rect 4973 -757 5019 -715
rect 4885 -856 4931 -757
rect 5061 -769 5089 -715
rect 5123 -721 5177 -715
rect 5149 -757 5177 -721
rect 4970 -779 5022 -773
rect 4970 -837 5022 -831
rect 4735 -928 4787 -925
rect 4735 -931 4849 -928
rect 4787 -940 4849 -931
rect 4787 -974 4805 -940
rect 4839 -974 4849 -940
rect 4903 -943 4931 -856
rect 5142 -940 5201 -928
rect 4903 -971 5107 -943
rect 4787 -983 4849 -974
rect 4735 -986 4849 -983
rect 4735 -989 4787 -986
rect 4970 -1084 5022 -1078
rect 4970 -1142 5022 -1136
rect 4815 -1195 4843 -1158
rect 4815 -1201 4875 -1195
rect 4903 -1201 4931 -1156
rect 4973 -1201 5019 -1158
rect 4815 -1235 4829 -1201
rect 4863 -1235 5019 -1201
rect 5079 -1185 5107 -971
rect 5142 -974 5154 -940
rect 5188 -974 5201 -940
rect 5142 -986 5201 -974
rect 5149 -1185 5177 -1119
rect 5079 -1201 5177 -1185
rect 5079 -1213 5129 -1201
rect 4815 -1241 5019 -1235
rect 4973 -1319 5019 -1241
rect 5121 -1235 5129 -1213
rect 5163 -1213 5177 -1201
rect 5163 -1235 5169 -1213
rect 5121 -1247 5169 -1235
rect 4735 -1491 4787 -1485
rect 4815 -1497 4843 -1419
rect 4885 -1497 4913 -1419
rect 5061 -1497 5089 -1419
rect 5149 -1497 5177 -1419
rect 5205 -1491 5257 -1485
rect 4787 -1503 4913 -1497
rect 4787 -1526 4829 -1503
rect 4815 -1537 4829 -1526
rect 4863 -1526 4913 -1503
rect 4941 -1503 5205 -1497
rect 4863 -1537 4875 -1526
rect 4815 -1543 4875 -1537
rect 4941 -1537 4953 -1503
rect 4987 -1525 5129 -1503
rect 4987 -1537 4999 -1525
rect 4941 -1543 4999 -1537
rect 5117 -1537 5129 -1525
rect 5163 -1525 5205 -1503
rect 5163 -1537 5177 -1525
rect 5117 -1543 5177 -1537
rect 4735 -1549 4787 -1543
rect 5205 -1549 5257 -1543
<< via1 >>
rect 4994 -379 5046 -377
rect 4994 -413 5005 -379
rect 5005 -413 5039 -379
rect 5039 -413 5046 -379
rect 4994 -429 5046 -413
rect 5058 -575 5110 -523
rect 4970 -831 5022 -779
rect 4735 -983 4787 -931
rect 4970 -1136 5022 -1084
rect 4735 -1543 4787 -1491
rect 5205 -1543 5257 -1491
<< metal2 >>
rect 4994 -371 5047 -363
rect 4994 -377 5257 -371
rect 5046 -429 5257 -377
rect 4994 -435 5046 -429
rect 5058 -523 5110 -517
rect 5058 -608 5110 -575
rect 4735 -660 5110 -608
rect 4735 -931 4787 -660
rect 4735 -1491 4787 -983
rect 4970 -779 5022 -773
rect 4970 -1084 5022 -831
rect 4970 -1142 5022 -1136
rect 4735 -1549 4787 -1543
rect 5205 -1491 5257 -429
rect 5205 -1549 5257 -1543
use sky130_fd_pr__nfet_01v8_6J3TAM  sky130_fd_pr__nfet_01v8_6J3TAM_0
timestamp 1730478237
transform 1 0 5128 0 1 -807
box -73 -76 73 76
use sky130_fd_pr__nfet_01v8_6J3TAM  sky130_fd_pr__nfet_01v8_6J3TAM_1
timestamp 1730478237
transform 1 0 4952 0 1 -547
box -73 -76 73 76
use sky130_fd_pr__nfet_01v8_6J3TAM  sky130_fd_pr__nfet_01v8_6J3TAM_2
timestamp 1730478237
transform 1 0 5040 0 1 -547
box -73 -76 73 76
use sky130_fd_pr__nfet_01v8_6J3TAM  sky130_fd_pr__nfet_01v8_6J3TAM_3
timestamp 1730478237
transform 1 0 4864 0 1 -547
box -73 -76 73 76
use sky130_fd_pr__nfet_01v8_6J3TAM  sky130_fd_pr__nfet_01v8_6J3TAM_4
timestamp 1730478237
transform 1 0 5128 0 1 -1109
box -73 -76 73 76
use sky130_fd_pr__nfet_01v8_6J3TAM  sky130_fd_pr__nfet_01v8_6J3TAM_5
timestamp 1730478237
transform 1 0 4952 0 1 -807
box -73 -76 73 76
use sky130_fd_pr__nfet_01v8_6J3TAM  sky130_fd_pr__nfet_01v8_6J3TAM_6
timestamp 1730478237
transform 1 0 5040 0 1 -807
box -73 -76 73 76
use sky130_fd_pr__nfet_01v8_6J3TAM  sky130_fd_pr__nfet_01v8_6J3TAM_7
timestamp 1730478237
transform 1 0 4864 0 1 -807
box -73 -76 73 76
use sky130_fd_pr__nfet_01v8_6J3TAM  sky130_fd_pr__nfet_01v8_6J3TAM_8
timestamp 1730478237
transform 1 0 4864 0 1 -1109
box -73 -76 73 76
use sky130_fd_pr__nfet_01v8_6J3TAM  sky130_fd_pr__nfet_01v8_6J3TAM_9
timestamp 1730478237
transform 1 0 4952 0 1 -1109
box -73 -76 73 76
use sky130_fd_pr__nfet_01v8_6J3TAM  sky130_fd_pr__nfet_01v8_6J3TAM_10
timestamp 1730478237
transform 1 0 5040 0 1 -1109
box -73 -76 73 76
use sky130_fd_pr__nfet_01v8_6J3TAM  sky130_fd_pr__nfet_01v8_6J3TAM_11
timestamp 1730478237
transform 1 0 5128 0 1 -547
box -73 -76 73 76
use sky130_fd_pr__nfet_01v8_6J3TAM  sky130_fd_pr__nfet_01v8_6J3TAM_12
timestamp 1730478237
transform -1 0 4952 0 -1 -1369
box -73 -76 73 76
use sky130_fd_pr__nfet_01v8_6J3TAM  sky130_fd_pr__nfet_01v8_6J3TAM_13
timestamp 1730478237
transform -1 0 5040 0 -1 -1369
box -73 -76 73 76
use sky130_fd_pr__nfet_01v8_6J3TAM  sky130_fd_pr__nfet_01v8_6J3TAM_14
timestamp 1730478237
transform -1 0 5128 0 -1 -1369
box -73 -76 73 76
use sky130_fd_pr__nfet_01v8_6J3TAM  sky130_fd_pr__nfet_01v8_6J3TAM_15
timestamp 1730478237
transform -1 0 4864 0 -1 -1369
box -73 -76 73 76
<< labels >>
flabel metal2 s 4996 -1018 4996 -1018 0 FreeSans 320 0 0 0 VDDA
port 1 nsew
flabel locali s 4997 -313 4997 -313 0 FreeSans 320 0 0 0 VSSA
port 5 nsew
flabel metal1 s 4846 -699 4846 -699 0 FreeSans 320 0 0 0 VPBT3
port 4 nsew
flabel metal2 s 4761 -1018 4761 -1018 0 FreeSans 320 0 0 0 VPBT1
port 2 nsew
flabel metal2 s 5232 -1018 5232 -1018 0 FreeSans 320 0 0 0 VPBT2
port 3 nsew
<< end >>
