magic
tech sky130A
timestamp 1730569521
<< nmos >>
rect -15 -25 15 25
<< ndiff >>
rect -44 19 -15 25
rect -44 -19 -38 19
rect -21 -19 -15 19
rect -44 -25 -15 -19
rect 15 19 44 25
rect 15 -19 21 19
rect 38 -19 44 19
rect 15 -25 44 -19
<< ndiffc >>
rect -38 -19 -21 19
rect 21 -19 38 19
<< poly >>
rect -15 25 15 38
rect -15 -38 15 -25
<< locali >>
rect -38 19 -21 27
rect -38 -27 -21 -19
rect 21 19 38 27
rect 21 -27 38 -19
<< viali >>
rect -38 -19 -21 19
rect 21 -19 38 19
<< metal1 >>
rect -41 19 -18 25
rect -41 -19 -38 19
rect -21 -19 -18 19
rect -41 -25 -18 -19
rect 18 19 41 25
rect 18 -19 21 19
rect 38 -19 41 19
rect 18 -25 41 -19
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
