magic
tech sky130A
magscale 1 2
timestamp 1730780526
<< nwell >>
rect 1301 216 1439 262
<< pwell >>
rect 3795 809 3991 875
<< locali >>
rect 1561 2225 1757 2291
rect 3795 809 3991 875
<< viali >>
rect 4205 2768 4239 2866
rect 3431 428 3625 530
rect 1313 234 1347 332
<< metal1 >>
rect 1277 3102 1678 3258
rect 1730 3102 3906 3258
rect 3958 3102 4275 3258
rect 621 3022 627 3074
rect 679 3022 1932 3074
rect 4239 2918 4870 2970
rect 4922 2918 4928 2970
rect 4129 2866 4251 2884
rect 4129 2838 4205 2866
rect 4193 2768 4205 2838
rect 4239 2768 4251 2866
rect 4193 2761 4251 2768
rect 1672 2232 1678 2284
rect 3795 861 3875 875
rect 3795 809 3817 861
rect 3869 809 3875 861
rect 3419 530 3637 536
rect 3419 428 3431 530
rect 3625 428 3637 530
rect 3419 422 3637 428
rect 1301 332 1359 339
rect 1301 234 1313 332
rect 1347 262 1359 332
rect 1347 234 1439 262
rect 1301 216 1439 234
rect 1575 130 4870 182
rect 4922 130 4928 182
rect 1277 -158 3431 -2
rect 3625 -158 4275 -2
<< via1 >>
rect 1678 3102 1730 3258
rect 3906 3102 3958 3258
rect 627 3022 679 3074
rect 4870 2918 4922 2970
rect 1678 2232 1730 2284
rect 3817 809 3869 861
rect 3431 428 3625 530
rect 4870 130 4922 182
rect 3431 -158 3625 -2
<< metal2 >>
rect 1678 3258 1730 3264
rect 627 3074 679 3080
rect 627 91 679 3022
rect 1678 2284 1730 3102
rect 3906 3258 3958 3264
rect 3906 2702 3958 3102
rect 4870 2970 4922 2976
rect 1678 1866 1730 2232
rect 1594 1814 1730 1866
rect 1594 1425 1646 1814
rect 3906 1283 3958 1669
rect 3817 1231 3958 1283
rect 3817 861 3869 1231
rect 3817 803 3869 809
rect 557 17 679 91
rect 3431 530 3625 536
rect 3431 -2 3625 428
rect 4870 182 4922 2918
rect 4870 124 4922 130
rect 3431 -164 3625 -158
use sh_bsw3  sh_bsw3_0 ~/sky130_projects/UNIC-CASS-2024/magic
timestamp 1730778869
transform -1 0 4275 0 -1 2708
box -1280 -375 2998 1604
use sh_bsw3  sh_bsw3_1
timestamp 1730778869
transform 1 0 1277 0 1 392
box -1280 -375 2998 1604
<< labels >>
flabel metal1 s 1277 3178 1277 3178 3 FreeSans 480 0 0 0 VDDA
port 1 e
flabel metal1 s 1113 153 1113 153 3 FreeSans 480 0 0 0 CLKS
port 2 e
flabel metal1 s 545 50 545 50 3 FreeSans 480 0 0 0 CLKSB
port 3 e
flabel metal1 s 2626 2850 2626 2850 3 FreeSans 480 0 0 0 VIP
port 4 e
flabel metal1 s 2626 249 2626 249 3 FreeSans 480 0 0 0 VIN
port 5 e
flabel metal1 s 1277 -86 1277 -86 3 FreeSans 480 0 0 0 VSSA
port 6 e
flabel metal2 s 2776 2956 2776 2956 3 FreeSans 480 0 0 0 VCP
port 7 e
flabel metal2 s 2775 144 2775 144 3 FreeSans 480 0 0 0 VCN
port 8 e
<< end >>
