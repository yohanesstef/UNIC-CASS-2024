magic
tech sky130A
magscale 1 2
timestamp 1730800306
<< nwell >>
rect 1003 1003 1055 1067
rect 918 957 964 985
rect 1094 929 1140 985
<< pwell >>
rect 1372 861 1626 1455
rect 686 791 2316 861
rect 536 776 2316 791
rect 536 770 2338 776
rect 536 740 1982 770
rect 600 0 1982 740
rect 2068 0 2338 770
rect 2629 85 2681 134
<< pdiff >>
rect 1045 1009 1055 1036
<< viali >>
rect 1262 387 1333 421
rect 1673 355 1744 389
<< metal1 >>
rect -196 1342 -183 1436
rect -131 1342 635 1436
rect 739 1342 745 1436
rect 1003 1303 1055 1309
rect 1003 1245 1055 1251
rect 766 1132 772 1184
rect 824 1132 1066 1184
rect 1003 1061 1055 1067
rect 1003 1003 1055 1009
rect 918 957 964 985
rect 1094 957 1140 985
rect -39 917 138 919
rect -39 825 -31 917
rect 25 825 138 917
rect 918 901 1140 957
rect -39 819 138 825
rect 2392 806 2450 811
rect 1003 791 1055 797
rect -756 690 -750 742
rect -694 690 196 742
rect 536 687 1003 791
rect 1003 681 1055 687
rect 1091 791 1143 797
rect 2392 791 2456 806
rect 1143 687 1271 791
rect 1323 687 1682 791
rect 1734 762 2456 791
rect 1734 687 2398 762
rect 2450 687 2456 762
rect 1091 681 1143 687
rect 879 595 885 647
rect 937 644 943 647
rect 2233 644 2239 647
rect 937 598 2239 644
rect 937 595 943 598
rect 2233 595 2239 598
rect 2291 595 2297 647
rect -40 386 -34 438
rect 18 386 552 438
rect 604 386 610 438
rect 766 382 772 434
rect 824 382 1024 434
rect 1265 427 1271 431
rect 1250 421 1271 427
rect 1323 427 1329 431
rect 1323 421 1345 427
rect 1250 387 1262 421
rect 1333 387 1345 421
rect 1250 381 1271 387
rect 1265 379 1271 381
rect 1323 381 1345 387
rect 1667 398 1750 401
rect 1667 389 1682 398
rect 1734 389 1750 398
rect 1323 379 1329 381
rect 1667 355 1673 389
rect 1744 355 1750 389
rect 1667 346 1682 355
rect 1734 346 1750 355
rect 1667 343 1750 346
rect 1996 287 2048 293
rect 1996 229 2048 235
rect 2635 134 2681 183
rect 629 50 635 102
rect 739 50 1181 102
rect 1233 50 1765 102
rect 1817 50 1823 102
rect 2233 44 2239 96
rect 2291 93 2297 96
rect 2629 93 2681 134
rect 2291 47 2681 93
rect 2291 44 2297 47
rect 766 -42 772 -36
rect 158 -88 772 -42
rect 824 -88 1996 -36
rect 2048 -88 2054 -36
rect 229 -176 235 -124
rect 287 -176 293 -124
rect 360 -210 418 -118
rect 454 -182 635 -130
rect 739 -182 745 -130
rect 1349 -168 1355 -116
rect 1407 -168 1591 -116
rect 1643 -168 1649 -116
rect -164 -262 -158 -210
rect -102 -262 418 -210
rect -889 -366 -880 -314
rect -824 -366 885 -314
rect 937 -366 943 -314
<< via1 >>
rect -183 1342 -131 1436
rect 635 1342 739 1436
rect 1003 1251 1055 1303
rect 772 1132 824 1184
rect 1003 1009 1055 1061
rect -31 825 25 917
rect -750 690 -694 742
rect 1003 687 1055 791
rect 1091 687 1143 791
rect 1271 687 1323 791
rect 1682 687 1734 791
rect 2398 687 2450 762
rect 885 595 937 647
rect 2239 595 2291 647
rect -34 386 18 438
rect 552 386 604 438
rect 772 382 824 434
rect 1271 421 1323 431
rect 1271 387 1323 421
rect 1271 379 1323 387
rect 1682 389 1734 398
rect 1682 355 1734 389
rect 1682 346 1734 355
rect 1996 235 2048 287
rect 635 50 739 102
rect 1181 50 1233 102
rect 1765 50 1817 102
rect 2239 44 2291 96
rect 772 -88 824 -36
rect 1996 -88 2048 -36
rect 235 -176 287 -124
rect 635 -182 739 -130
rect 1355 -168 1407 -116
rect 1591 -168 1643 -116
rect -158 -262 -102 -210
rect -880 -366 -824 -314
rect 885 -366 937 -314
<< metal2 >>
rect -196 1570 -127 1579
rect -196 1498 -189 1570
rect -133 1498 -127 1570
rect -196 1436 -127 1498
rect -196 1342 -183 1436
rect -131 1342 -127 1436
rect -196 1333 -127 1342
rect 635 1436 739 1442
rect -31 1214 25 1223
rect -31 917 25 1097
rect -31 819 25 825
rect -750 742 -694 748
rect -750 203 -694 690
rect -750 77 -694 86
rect -34 438 18 444
rect -34 210 18 386
rect -34 201 25 210
rect -34 84 -31 201
rect -34 79 25 84
rect -31 75 25 79
rect 317 -124 369 404
rect 552 160 604 288
rect 201 -176 235 -124
rect 287 -176 369 -124
rect 635 102 739 1342
rect 1003 1303 1055 1309
rect 635 -130 739 50
rect 772 1184 824 1190
rect 772 434 824 1132
rect 1003 1061 1055 1251
rect 1003 791 1055 1009
rect 1003 681 1055 687
rect 1091 791 1143 1139
rect 1091 681 1143 687
rect 1271 791 1323 797
rect 772 -36 824 382
rect 772 -94 824 -88
rect 885 647 937 654
rect 635 -188 739 -182
rect -158 -206 -95 -197
rect -158 -210 -151 -206
rect -163 -262 -158 -210
rect -163 -271 -95 -262
rect -880 -310 -824 -301
rect -880 -375 -824 -366
rect 885 -314 937 595
rect 1271 431 1323 687
rect 1271 373 1323 379
rect 1682 791 1734 797
rect 1682 398 1734 687
rect 2239 647 2291 653
rect 2239 589 2291 595
rect 1181 102 1233 234
rect 1181 44 1233 50
rect 1355 -116 1407 377
rect 1355 -174 1407 -168
rect 1473 -228 1525 373
rect 1591 -116 1643 360
rect 1682 340 1734 346
rect 1765 102 1817 343
rect 1765 44 1817 50
rect 1996 287 2048 293
rect 1996 -36 2048 235
rect 2242 102 2288 589
rect 2239 96 2291 102
rect 2239 38 2291 44
rect 1996 -94 2048 -88
rect 1591 -174 1643 -168
rect 885 -372 937 -366
<< via2 >>
rect -189 1498 -133 1570
rect -31 1097 25 1214
rect -750 86 -694 203
rect -31 84 25 201
rect -151 -210 -95 -206
rect -151 -262 -102 -210
rect -102 -262 -95 -210
rect -880 -314 -824 -310
rect -880 -366 -824 -314
<< metal3 >>
rect -196 1570 -127 1579
rect -196 1498 -189 1570
rect -133 1498 -127 1570
rect -40 1214 31 1226
rect -40 1097 -39 1214
rect 25 1097 31 1214
rect -40 1085 31 1097
rect -758 203 -687 214
rect -694 86 -687 203
rect -758 73 -687 86
rect -40 201 31 212
rect 25 84 31 201
rect -40 71 31 84
rect -880 -305 -820 10
rect -160 -201 -100 0
rect -160 -206 -90 -201
rect -160 -262 -151 -206
rect -95 -262 -90 -206
rect -160 -271 -90 -262
rect -886 -310 -816 -305
rect -886 -366 -880 -310
rect -824 -366 -816 -310
rect -886 -376 -816 -366
<< via3 >>
rect -39 1097 -31 1214
rect -31 1097 25 1214
rect -758 86 -750 203
rect -750 86 -694 203
rect -40 84 -31 201
rect -31 84 24 201
<< metal4 >>
rect -179 1214 31 1219
rect -179 1097 -39 1214
rect 25 1097 31 1214
rect -179 1091 31 1097
rect -1073 273 -1069 401
rect -758 207 -687 214
rect -957 203 -687 207
rect -957 86 -758 203
rect -694 86 -687 203
rect -957 79 -687 86
rect -179 201 25 207
rect -179 84 -40 201
rect 24 84 25 201
rect -179 79 25 84
rect -758 73 -687 79
use cap_bsw  cap_bsw_1
timestamp 1730798039
transform 0 -1 -1234 1 0 -1462
box 1462 -1134 3246 66
use inv_bsw  inv_bsw_0
timestamp 1730718786
transform 0 -1 563 1 0 -215
box -3 -123 215 563
use ncell_bsw  ncell_bsw_1
timestamp 1730778869
transform 1 0 -4653 0 1 1676
box 4653 -1676 5339 -261
use ncell_bsw_dischrg  ncell_bsw_dischrg_0
timestamp 1730741927
transform 1 0 2450 0 1 1725
box -138 -1725 548 -824
use ncell_bsw_sw  ncell_bsw_sw_1
timestamp 1730741762
transform 1 0 1311 0 1 3662
box -503 -3662 879 -2886
use pcell_bsw_dischrg  pcell_bsw_dischrg_0
timestamp 1730722715
transform 1 0 75 0 1 1310
box 611 -449 1297 145
<< labels >>
flabel metal2 s 342 -3 342 -3 0 FreeSans 320 0 0 0 VDDA
port 1 nsew
flabel metal1 s 162 -237 162 -237 0 FreeSans 320 0 0 0 CLKS
port 2 nsew
flabel metal1 s 161 -342 161 -342 0 FreeSans 320 0 0 0 CLKSB
port 3 nsew
flabel metal2 s 1381 -23 1381 -23 0 FreeSans 320 0 0 0 VI
port 4 nsew
flabel locali s 570 54 570 54 0 FreeSans 320 0 0 0 VSSA
port 5 nsew
flabel metal2 s 1499 -215 1499 -215 0 FreeSans 320 0 0 0 VO
port 6 nsew
<< end >>
