magic
tech sky130A
magscale 1 2
timestamp 1729091911
<< pwell >>
rect 3264 -84 3333 -13
rect 2402 -322 2504 -127
rect 3318 -375 3370 -254
rect 3824 -332 4824 -280
<< locali >>
rect -616 1556 5197 1576
rect -616 1496 -596 1556
rect 5177 1496 5197 1556
rect -616 1377 5197 1496
rect -616 1307 856 1377
rect -616 827 -382 1307
rect 532 827 856 1307
rect 891 829 1047 1229
rect -616 609 856 827
rect 1278 609 5197 1377
rect -616 481 5197 609
rect -616 18 5197 280
rect -616 -98 768 18
rect -616 -400 -382 -98
rect 532 -400 768 -98
rect 1050 -98 3156 18
rect 1050 -400 1172 -98
rect 3034 -400 3156 -98
rect 3438 -88 5197 18
rect 3438 -400 3684 -88
rect 4902 -400 5197 -88
rect -616 -520 5197 -400
rect -616 -580 -596 -520
rect 5177 -580 5197 -520
rect -616 -600 5197 -580
<< viali >>
rect -596 1496 5177 1556
rect -596 -580 5177 -520
<< metal1 >>
rect -616 1556 5197 1576
rect -616 1496 -596 1556
rect 5177 1496 5197 1556
rect -616 1476 5197 1496
rect -308 1229 -262 1476
rect 8 1229 54 1476
rect -174 977 -100 1229
rect 96 977 216 1229
rect 324 1210 370 1476
rect 458 977 532 1229
rect -168 930 -100 977
rect 148 936 216 977
rect -274 463 -208 929
rect -617 311 -208 463
rect -274 -200 -208 311
rect -168 880 108 930
rect -168 118 -100 880
rect -168 33 -161 118
rect -108 33 -100 118
rect -168 -150 -100 33
rect 42 -150 108 880
rect -168 -200 108 -150
rect 148 880 424 936
rect 148 598 216 880
rect 148 407 155 598
rect 210 407 216 598
rect 148 -150 216 407
rect 358 -150 424 880
rect 148 -200 424 -150
rect 464 782 532 977
rect 464 697 471 782
rect 524 697 532 782
rect -168 -238 -100 -200
rect 148 -238 216 -200
rect 464 -238 532 697
rect 836 829 1047 1229
rect 1084 932 1137 938
rect 1084 841 1137 847
rect 836 -60 888 829
rect 1034 784 1100 788
rect 1028 732 1034 784
rect 1100 732 1106 784
rect 1169 -60 1292 1476
rect -308 -500 -262 -238
rect -220 -322 -100 -238
rect 8 -500 54 -238
rect 96 -322 216 -238
rect 412 -322 532 -238
rect 590 -61 888 -60
rect 590 -259 612 -61
rect 772 -259 888 -61
rect 590 -260 888 -259
rect 930 -260 1292 -60
rect 1334 1221 1453 1224
rect 1334 1014 1344 1221
rect 1447 1014 1453 1221
rect 1334 -176 1453 1014
rect 1485 -60 1608 1476
rect 2402 846 2429 931
rect 2482 846 2503 931
rect 2120 699 2127 784
rect 2180 699 2187 784
rect 1333 -260 1488 -176
rect 1524 -260 1608 -60
rect 1710 357 1804 363
rect 1710 178 1722 357
rect 1793 178 1804 357
rect 1710 -176 1804 178
rect 1650 -260 1804 -176
rect 1912 119 1978 124
rect 1912 34 1918 119
rect 1971 34 1978 119
rect 1912 -200 1978 34
rect 2120 -238 2187 699
rect 2402 425 2503 846
rect 2402 -29 2504 425
rect 2396 -35 2504 -29
rect 2396 -93 2402 -35
rect 2454 -93 2504 -35
rect 2396 -99 2504 -93
rect 2402 -150 2504 -99
rect 2228 -200 2504 -150
rect 2544 -200 2610 1476
rect 2860 118 2926 126
rect 2860 33 2867 118
rect 2920 33 2926 118
rect 2860 -200 2926 33
rect 3264 -19 3792 -13
rect 3264 -77 3273 -19
rect 3325 -77 3792 -19
rect 3264 -84 3792 -77
rect 2402 -238 2504 -200
rect 1454 -298 1488 -260
rect 324 -399 370 -322
rect 876 -370 1346 -298
rect 1454 -338 1662 -298
rect 1710 -370 1804 -260
rect 316 -405 380 -399
rect 876 -400 1804 -370
rect 1872 -393 1924 -238
rect 1866 -399 1930 -393
rect 316 -463 322 -405
rect 374 -463 380 -405
rect 1866 -457 1872 -399
rect 1924 -457 1930 -399
rect 1866 -463 1930 -457
rect 316 -469 380 -463
rect 1966 -500 2018 -238
rect 2120 -322 2240 -238
rect 2284 -337 2348 -238
rect 2402 -322 2556 -238
rect 2597 -322 2870 -237
rect 2284 -395 2290 -337
rect 2342 -395 2348 -337
rect 2284 -401 2348 -395
rect 2914 -500 2960 -238
rect 3222 -331 3276 -122
rect 3211 -337 3276 -331
rect 3211 -395 3217 -337
rect 3269 -395 3276 -337
rect 3211 -401 3276 -395
rect 3318 -323 3370 -122
rect 3684 -277 3792 -84
rect 3823 -207 5197 -54
rect 3824 -208 5197 -207
rect 3824 -323 4824 -280
rect 3318 -332 4824 -323
rect 3318 -434 5197 -332
rect -616 -520 5197 -500
rect -616 -580 -596 -520
rect 5177 -580 5197 -520
rect -616 -600 5197 -580
<< via1 >>
rect -161 33 -108 118
rect 155 407 210 598
rect 471 697 524 782
rect 1084 847 1137 932
rect 1034 732 1100 784
rect 612 -259 772 -61
rect 1344 1014 1447 1221
rect 2429 846 2482 931
rect 2127 699 2180 784
rect 1722 178 1793 357
rect 1918 34 1971 119
rect 2402 -93 2454 -35
rect 2867 33 2920 118
rect 3273 -77 3325 -19
rect 322 -463 374 -405
rect 1872 -457 1924 -399
rect 2290 -395 2342 -337
rect 3217 -395 3269 -337
<< metal2 >>
rect 1335 1221 2424 1226
rect 1335 1014 1344 1221
rect 1447 1210 2424 1221
rect 1447 1019 2289 1210
rect 2419 1019 2424 1210
rect 1447 1014 2424 1019
rect 1335 1007 2424 1014
rect 1084 932 2503 938
rect 1137 931 2503 932
rect 1137 847 2429 931
rect 1084 846 2429 847
rect 2482 846 2503 931
rect 1084 841 2503 846
rect 464 782 1034 784
rect 464 697 471 782
rect 524 732 1034 782
rect 1100 732 2127 784
rect 524 699 2127 732
rect 2180 699 2187 784
rect 524 697 2187 699
rect 464 693 2187 697
rect 147 407 155 598
rect 210 407 2657 598
rect 1710 357 2237 363
rect 1710 178 1722 357
rect 1793 178 2237 357
rect 1710 172 2237 178
rect 2367 172 2392 363
rect 2542 302 2657 407
rect 2542 288 4003 302
rect 2542 224 2549 288
rect 3987 224 4003 288
rect 2542 212 4003 224
rect -168 119 2926 124
rect -168 118 1918 119
rect -168 33 -161 118
rect -108 111 1918 118
rect 1971 118 2926 119
rect 1971 111 2867 118
rect -108 47 637 111
rect 2075 47 2867 111
rect -108 34 1918 47
rect 1971 34 2867 47
rect -108 33 2867 34
rect 2920 33 2926 118
rect -168 27 2926 33
rect 3264 -19 3333 -13
rect 3264 -29 3273 -19
rect 2396 -35 3273 -29
rect 600 -259 612 -61
rect 772 -259 781 -61
rect 2396 -93 2402 -35
rect 2454 -77 3273 -35
rect 3325 -77 3333 -19
rect 2454 -93 3333 -77
rect 2396 -99 3333 -93
rect 2282 -337 3276 -331
rect 22 -405 391 -398
rect 1866 -399 1930 -393
rect 1866 -405 1872 -399
rect 22 -463 322 -405
rect 374 -457 1872 -405
rect 1924 -405 1930 -399
rect 2282 -395 2290 -337
rect 2342 -395 3217 -337
rect 3269 -395 3276 -337
rect 2282 -401 3276 -395
rect 2282 -405 2349 -401
rect 1924 -457 2349 -405
rect 374 -463 2349 -457
rect 22 -475 2349 -463
rect 22 -625 391 -475
rect 22 -665 37 -625
rect 21 -800 37 -665
rect 102 -800 391 -625
rect 21 -814 391 -800
<< via2 >>
rect 2289 1019 2419 1210
rect 2237 172 2367 363
rect 2549 224 3987 288
rect 637 47 1918 111
rect 1918 47 1971 111
rect 1971 47 2075 111
rect 612 -259 772 -61
rect 37 -800 102 -625
<< metal3 >>
rect 2283 1210 2424 1227
rect 2283 1019 2289 1210
rect 2419 1019 2424 1210
rect 2283 1008 2424 1019
rect 2231 605 2374 624
rect 2231 414 2238 605
rect 2368 414 2374 605
rect 2231 363 2374 414
rect 2231 172 2237 363
rect 2367 172 2374 363
rect 2231 164 2374 172
rect 606 -61 778 -54
rect 606 -259 612 -61
rect 772 -259 778 -61
rect 606 -265 778 -259
<< via3 >>
rect 2289 1019 2419 1210
rect 2238 414 2368 605
rect 612 -259 772 -61
<< metal4 >>
rect 2283 1210 2641 1227
rect 2283 1019 2289 1210
rect 2419 1019 2641 1210
rect 2283 1008 2641 1019
rect 1974 605 2375 624
rect 1974 414 2238 605
rect 2368 414 2375 605
rect 1974 398 2375 414
rect 552 -61 835 -60
rect 552 -259 612 -61
rect 772 -259 835 -61
rect 552 -713 835 -259
use sky130_fd_pr__nfet_01v8_L78EGD  sky130_fd_pr__nfet_01v8_L78EGD_0
timestamp 1729068740
transform 1 0 -241 0 1 -249
box -211 -221 211 221
use sky130_fd_pr__nfet_01v8_TK2CNP  sky130_fd_pr__nfet_01v8_TK2CNP_0
timestamp 1729087186
transform 0 -1 4293 1 0 -244
box -226 -679 226 679
use sky130_fd_pr__pfet_01v8_LCNWMQ  sky130_fd_pr__pfet_01v8_LCNWMQ_0
timestamp 1729068740
transform 1 0 391 0 1 1067
box -211 -310 211 310
use sky130_fd_pr__cap_mim_m3_1_5XYVA6  XC1
timestamp 1729087186
transform 0 1 1356 -1 0 920
box -893 -747 893 747
use sky130_fd_pr__cap_mim_m3_1_5XY9G7  XC2
timestamp 1729068740
transform 0 1 3271 -1 0 921
box -893 -747 893 747
use sky130_fd_pr__cap_mim_m3_1_QEFW4K  XC3
timestamp 1729068740
transform -1 0 2435 0 -1 -2874
box -2417 -2271 2417 2271
use sky130_fd_pr__nfet_01v8_L78EGD  XM1
timestamp 1729068740
transform -1 0 1313 0 -1 -249
box -211 -221 211 221
use sky130_fd_pr__pfet_01v8_M4BBJH  XM2
timestamp 1729068740
transform 1 0 1067 0 1 993
box -211 -384 211 384
use sky130_fd_pr__nfet_01v8_L78EGD  XM3
timestamp 1729068740
transform -1 0 1629 0 -1 -249
box -211 -221 211 221
use sky130_fd_pr__nfet_01v8_7XY3PK  XM4
timestamp 1729068740
transform -1 0 909 0 -1 -191
box -211 -279 211 279
use sky130_fd_pr__nfet_01v8_L78EGD  XM5
timestamp 1729068740
transform 1 0 1945 0 1 -249
box -211 -221 211 221
use sky130_fd_pr__nfet_01v8_L78EGD  XM7
timestamp 1729068740
transform 1 0 391 0 1 -249
box -211 -221 211 221
use sky130_fd_pr__nfet_01v8_L78EGD  XM8
timestamp 1729068740
transform 1 0 2577 0 1 -249
box -211 -221 211 221
use sky130_fd_pr__nfet_01v8_L78EGD  XM9
timestamp 1729068740
transform 1 0 2893 0 1 -249
box -211 -221 211 221
use sky130_fd_pr__nfet_01v8_L78EGD  XM10
timestamp 1729068740
transform 1 0 2261 0 1 -249
box -211 -221 211 221
use sky130_fd_pr__nfet_01v8_7XY3PK  XM11
timestamp 1729068740
transform 1 0 3297 0 1 -191
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_LCNWMQ  XM13
timestamp 1729068740
transform 1 0 -241 0 1 1067
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_LCNWMQ  XM15
timestamp 1729068740
transform 1 0 75 0 1 1067
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_L78EGD  XM16
timestamp 1729068740
transform 1 0 75 0 1 -249
box -211 -221 211 221
<< labels >>
flabel metal1 -617 382 -617 382 3 FreeSans 800 0 0 0 clk
port 1 e
flabel metal1 5197 -391 5197 -391 7 FreeSans 800 0 0 0 vdata
port 2 w
flabel metal1 -616 1524 -616 1524 3 FreeSans 800 0 0 0 VDD
port 3 e
flabel metal1 -616 -550 -616 -550 3 FreeSans 800 0 0 0 GND
port 4 e
flabel metal1 5197 -134 5197 -134 7 FreeSans 800 0 0 0 Vout
port 6 w
flabel metal1 s 3570 -50 3570 -50 0 FreeSans 800 0 0 0 vboot
<< end >>
