* NGSPICE file created from sh_bsw.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_275TTJ a_n15_n76# w_n109_n112# a_n73_n50# a_15_n50#
+ VSUBS
X0 a_15_n50# a_n15_n76# a_n73_n50# w_n109_n112# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
C0 w_n109_n112# a_n73_n50# 0.00578f
C1 a_n15_n76# a_15_n50# 0.003563f
C2 a_n15_n76# w_n109_n112# 0.022339f
C3 a_n15_n76# a_n73_n50# 0.003563f
C4 w_n109_n112# a_15_n50# 0.00578f
C5 a_n73_n50# a_15_n50# 0.082646f
C6 a_15_n50# VSUBS 0.070304f
C7 a_n73_n50# VSUBS 0.070304f
C8 a_n15_n76# VSUBS 0.043702f
C9 w_n109_n112# VSUBS 0.146496f
.ends

.subckt pcell_bsw_dischrg VPBT3 SWITCHING VBOOT VSUBS
Xsky130_fd_pr__pfet_01v8_275TTJ_6 VPBT3 VPBT3 VPBT3 VBOOT VSUBS sky130_fd_pr__pfet_01v8_275TTJ
Xsky130_fd_pr__pfet_01v8_275TTJ_7 SWITCHING VPBT3 VPBT3 VBOOT VSUBS sky130_fd_pr__pfet_01v8_275TTJ
Xsky130_fd_pr__pfet_01v8_275TTJ_0 SWITCHING VPBT3 VBOOT VPBT3 VSUBS sky130_fd_pr__pfet_01v8_275TTJ
Xsky130_fd_pr__pfet_01v8_275TTJ_1 SWITCHING VPBT3 VPBT3 VBOOT VSUBS sky130_fd_pr__pfet_01v8_275TTJ
Xsky130_fd_pr__pfet_01v8_275TTJ_3 VPBT3 VPBT3 VPBT3 VBOOT VSUBS sky130_fd_pr__pfet_01v8_275TTJ
Xsky130_fd_pr__pfet_01v8_275TTJ_2 SWITCHING VPBT3 VBOOT VPBT3 VSUBS sky130_fd_pr__pfet_01v8_275TTJ
Xsky130_fd_pr__pfet_01v8_275TTJ_4 VPBT3 VPBT3 VBOOT VPBT3 VSUBS sky130_fd_pr__pfet_01v8_275TTJ
Xsky130_fd_pr__pfet_01v8_275TTJ_5 VPBT3 VPBT3 VBOOT VPBT3 VSUBS sky130_fd_pr__pfet_01v8_275TTJ
C0 SWITCHING VBOOT 0.171013f
C1 VPBT3 VBOOT 0.283635f
C2 VPBT3 SWITCHING 0.293769f
C3 VBOOT VSUBS 0.169533f
C4 SWITCHING VSUBS 0.111275f
C5 VPBT3 VSUBS 2.478131f
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_VCTT89 m3_n386_n240# c1_n346_n200# VSUBS
X0 c1_n346_n200# m3_n386_n240# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
C0 m3_n386_n240# c1_n346_n200# 0.507132f
C1 c1_n346_n200# VSUBS 0.169673f
C2 m3_n386_n240# VSUBS 0.762748f
.ends

.subckt cap_bsw VPBT1 VNBT1 VPBT2 VPBT3 VNBT3 CLKS VSUBS
Xsky130_fd_pr__cap_mim_m3_1_VCTT89_0 VNBT3 VPBT3 VSUBS sky130_fd_pr__cap_mim_m3_1_VCTT89
Xsky130_fd_pr__cap_mim_m3_1_VCTT89_1 VNBT3 VPBT3 VSUBS sky130_fd_pr__cap_mim_m3_1_VCTT89
XXC1 VNBT1 VPBT1 VSUBS sky130_fd_pr__cap_mim_m3_1_VCTT89
XXC2 CLKS VPBT2 VSUBS sky130_fd_pr__cap_mim_m3_1_VCTT89
C0 CLKS VPBT1 0.012183f
C1 VNBT3 VPBT3 0.143473f
C2 VNBT1 CLKS 0.382401f
C3 VNBT1 VPBT3 0.13591f
C4 VNBT3 VNBT1 0.312674f
C5 VPBT1 VPBT2 0.084078f
C6 VNBT1 VPBT2 0.012183f
C7 CLKS VPBT3 0.13591f
C8 VNBT3 CLKS 0.312674f
C9 VPBT3 VSUBS 0.160558f
C10 VNBT3 VSUBS 1.011946f
C11 VPBT2 VSUBS 0.11587f
C12 CLKS VSUBS 0.424282f
C13 VPBT1 VSUBS 0.11587f
C14 VNBT1 VSUBS 0.424282f
.ends

.subckt sky130_fd_pr__nfet_01v8_QS6TK8 a_30_n50# a_n30_n76# a_n88_n50# VSUBS
X0 a_30_n50# a_n30_n76# a_n88_n50# VSUBS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.3
C0 a_n88_n50# a_30_n50# 0.061754f
C1 a_n30_n76# a_30_n50# 0.006618f
C2 a_n30_n76# a_n88_n50# 0.006618f
C3 a_30_n50# VSUBS 0.076817f
C4 a_n88_n50# VSUBS 0.076817f
C5 a_n30_n76# VSUBS 0.103343f
.ends

.subckt sky130_fd_pr__nfet_01v8_6J3TAM a_n15_n76# a_n73_n50# a_15_n50# VSUBS
X0 a_15_n50# a_n15_n76# a_n73_n50# VSUBS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
C0 a_n73_n50# a_15_n50# 0.082646f
C1 a_n15_n76# a_15_n50# 0.003563f
C2 a_n15_n76# a_n73_n50# 0.003563f
C3 a_15_n50# VSUBS 0.076084f
C4 a_n73_n50# VSUBS 0.076084f
C5 a_n15_n76# VSUBS 0.066041f
.ends

.subckt ncell_bsw_sw VI VBOOT VNBT1 VNBT3 SWITCHING VO VSSA
Xsky130_fd_pr__nfet_01v8_QS6TK8_0 VI VBOOT VNBT3 VSSA sky130_fd_pr__nfet_01v8_QS6TK8
Xsky130_fd_pr__nfet_01v8_QS6TK8_1 VO VBOOT VI VSSA sky130_fd_pr__nfet_01v8_QS6TK8
Xsky130_fd_pr__nfet_01v8_QS6TK8_2 VI VBOOT VO VSSA sky130_fd_pr__nfet_01v8_QS6TK8
Xsky130_fd_pr__nfet_01v8_QS6TK8_4 VI VI VI VSSA sky130_fd_pr__nfet_01v8_QS6TK8
Xsky130_fd_pr__nfet_01v8_QS6TK8_3 VNBT3 VBOOT VI VSSA sky130_fd_pr__nfet_01v8_QS6TK8
Xsky130_fd_pr__nfet_01v8_QS6TK8_5 VI VI VI VSSA sky130_fd_pr__nfet_01v8_QS6TK8
Xsky130_fd_pr__nfet_01v8_6J3TAM_10 SWITCHING SWITCHING SWITCHING VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_QS6TK8_6 VO VBOOT VI VSSA sky130_fd_pr__nfet_01v8_QS6TK8
Xsky130_fd_pr__nfet_01v8_QS6TK8_7 VI VBOOT VO VSSA sky130_fd_pr__nfet_01v8_QS6TK8
Xsky130_fd_pr__nfet_01v8_6J3TAM_0 VBOOT SWITCHING VNBT3 VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_1 VBOOT VNBT3 SWITCHING VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_2 VNBT1 VSSA VNBT3 VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_3 VNBT1 VNBT3 VSSA VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_4 VSSA VSSA VSSA VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_5 VSSA VSSA VSSA VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_6 SWITCHING SWITCHING SWITCHING VSSA sky130_fd_pr__nfet_01v8_6J3TAM
C0 VO VNBT3 0.002465f
C1 VNBT1 VNBT3 0.279574f
C2 SWITCHING VNBT3 0.076911f
C3 VO VI 0.327127f
C4 VBOOT VNBT3 0.3325f
C5 VNBT1 VI 0.29817f
C6 SWITCHING VI 0.007735f
C7 VBOOT VI 0.428361f
C8 VO VNBT1 0.002161f
C9 VO SWITCHING 0.001334f
C10 VO VBOOT 0.101863f
C11 SWITCHING VNBT1 0.894613f
C12 VBOOT VNBT1 0.090912f
C13 VBOOT SWITCHING 0.147106f
C14 VI VNBT3 0.533331f
C15 VNBT3 VSSA 0.497171f
C16 VI VSSA 0.528057f
C17 VNBT1 VSSA 0.862944f
C18 SWITCHING VSSA 1.479728f
C19 VBOOT VSSA 0.935003f
C20 VO VSSA 0.055615f
.ends

.subckt ncell_bsw_dischrg VDDA CLKSB VBOOT VSSA a_179_n1156#
Xsky130_fd_pr__nfet_01v8_6J3TAM_0 VBOOT VBOOT VBOOT VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_1 VSSA VSSA VSSA VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_2 CLKSB VSSA a_179_n1156# VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_3 VDDA a_179_n1156# VBOOT VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_4 VBOOT VBOOT VBOOT VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_5 VDDA VBOOT a_179_n1156# VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_6 CLKSB a_179_n1156# VSSA VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_7 VSSA VSSA VSSA VSSA sky130_fd_pr__nfet_01v8_6J3TAM
C0 CLKSB VSSA 0.053992f
C1 VDDA CLKSB 0.09168f
C2 CLKSB a_179_n1156# 0.135282f
C3 VDDA VSSA 0.030733f
C4 a_179_n1156# VSSA 0.003384f
C5 VDDA a_179_n1156# 0.08975f
C6 VBOOT CLKSB 0.335238f
C7 VBOOT VSSA 0.117288f
C8 VDDA VBOOT 0.105082f
C9 VBOOT a_179_n1156# 0.003556f
C10 VSSA 0 0.047349f
C11 a_179_n1156# 0 0.072735f
C12 CLKSB 0 0.601343f
C13 VBOOT 0 1.166181f
C14 VDDA 0 0.340207f
.ends

.subckt ncell_bsw VDDA VPBT1 VPBT2 VPBT3 VSSA
Xsky130_fd_pr__nfet_01v8_6J3TAM_10 VPBT1 VDDA VPBT3 VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_11 VPBT1 VPBT1 VPBT1 VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_12 VPBT2 VDDA VPBT1 VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_13 VPBT1 VPBT2 VDDA VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_14 VPBT2 VPBT2 VPBT2 VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_15 VPBT1 VPBT1 VPBT1 VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_0 VDDA VDDA VDDA VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_1 VPBT1 VPBT2 VDDA VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_2 VPBT2 VDDA VPBT1 VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_3 VPBT2 VPBT2 VPBT2 VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_4 VPBT3 VPBT3 VPBT3 VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_5 VPBT1 VPBT3 VDDA VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_6 VDDA VDDA VDDA VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_7 VPBT3 VPBT3 VPBT3 VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_8 VDDA VDDA VDDA VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_9 VDDA VDDA VDDA VSSA sky130_fd_pr__nfet_01v8_6J3TAM
C0 VPBT2 VDDA 0.222284f
C1 VPBT2 VPBT1 0.563039f
C2 VPBT3 VDDA 0.232497f
C3 VPBT1 VPBT3 0.336182f
C4 VPBT1 VDDA 0.596132f
C5 VPBT2 VPBT3 0.194492f
C6 VPBT3 VSSA 0.484194f
C7 VPBT1 VSSA 1.487454f
C8 VDDA VSSA 0.708267f
C9 VPBT2 VSSA 1.397263f
.ends

.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
C0 Y A 0.047605f
C1 VGND Y 0.099841f
C2 VPWR A 0.037031f
C3 VGND VPWR 0.033816f
C4 VPB A 0.045062f
C5 VGND VPB 0.009478f
C6 Y VPWR 0.127579f
C7 Y VPB 0.017744f
C8 VPWR VPB 0.054478f
C9 VGND A 0.040045f
C10 VGND VNB 0.251126f
C11 Y VNB 0.096099f
C12 VPWR VNB 0.218922f
C13 A VNB 0.166643f
C14 VPB VNB 0.338976f
.ends

.subckt sh_bsw VDDA CLKS CLKSB VI VSSA VO
Xpcell_bsw_dischrg_1 cap_bsw_1/VPBT3 ncell_bsw_sw_1/SWITCHING ncell_bsw_sw_1/VBOOT
+ VSSA pcell_bsw_dischrg
Xcap_bsw_1 cap_bsw_1/VPBT1 CLKSB cap_bsw_1/VPBT2 cap_bsw_1/VPBT3 cap_bsw_1/VNBT3 CLKS
+ VSSA cap_bsw
Xncell_bsw_sw_1 VI ncell_bsw_sw_1/VBOOT CLKSB cap_bsw_1/VNBT3 ncell_bsw_sw_1/SWITCHING
+ VO VSSA ncell_bsw_sw
Xncell_bsw_dischrg_1 VDDA CLKSB ncell_bsw_sw_1/VBOOT VSSA ncell_bsw_dischrg_1/a_179_n1156#
+ ncell_bsw_dischrg
Xncell_bsw_1 VDDA cap_bsw_1/VPBT1 cap_bsw_1/VPBT2 cap_bsw_1/VPBT3 VSSA ncell_bsw
Xsky130_fd_sc_hd__inv_1_0 CLKS cap_bsw_1/VNBT3 VSSA VDDA VDDA ncell_bsw_sw_1/SWITCHING
+ sky130_fd_sc_hd__inv_1
C0 cap_bsw_1/VPBT1 cap_bsw_1/VPBT2 1.122085f
C1 cap_bsw_1/VPBT1 cap_bsw_1/VNBT3 0.085121f
C2 cap_bsw_1/VPBT1 CLKS 0.124177f
C3 ncell_bsw_sw_1/VBOOT VI 0.078231f
C4 cap_bsw_1/VPBT3 ncell_bsw_sw_1/VBOOT 0.401711f
C5 VSSA VI 0.01058f
C6 cap_bsw_1/VPBT3 VSSA 0.665901f
C7 cap_bsw_1/VPBT1 VI 0.048922f
C8 cap_bsw_1/VPBT1 cap_bsw_1/VPBT3 0.046341f
C9 ncell_bsw_sw_1/VBOOT VO 0.003085f
C10 VDDA ncell_bsw_sw_1/SWITCHING 0.504446f
C11 ncell_bsw_sw_1/VBOOT CLKSB 0.10443f
C12 cap_bsw_1/VPBT2 ncell_bsw_sw_1/SWITCHING 0.084824f
C13 VSSA VO 0.006757f
C14 ncell_bsw_sw_1/SWITCHING cap_bsw_1/VNBT3 0.895623f
C15 CLKS ncell_bsw_sw_1/SWITCHING 0.688459f
C16 CLKSB VSSA 0.098445f
C17 ncell_bsw_dischrg_1/a_179_n1156# ncell_bsw_sw_1/SWITCHING 5.51e-20
C18 VDDA cap_bsw_1/VPBT2 0.304087f
C19 cap_bsw_1/VPBT1 VO 0.042758f
C20 VDDA cap_bsw_1/VNBT3 -0.006184f
C21 VDDA CLKS 0.060834f
C22 cap_bsw_1/VPBT1 CLKSB 0.457202f
C23 cap_bsw_1/VPBT2 cap_bsw_1/VNBT3 0.050391f
C24 CLKS cap_bsw_1/VPBT2 0.581513f
C25 VDDA ncell_bsw_dischrg_1/a_179_n1156# 4.71e-19
C26 CLKS cap_bsw_1/VNBT3 0.614317f
C27 ncell_bsw_dischrg_1/a_179_n1156# cap_bsw_1/VPBT2 2.66e-21
C28 ncell_bsw_dischrg_1/a_179_n1156# cap_bsw_1/VNBT3 0.006241f
C29 ncell_bsw_sw_1/SWITCHING VI 0.064143f
C30 cap_bsw_1/VPBT3 ncell_bsw_sw_1/SWITCHING 0.210561f
C31 VDDA VI 0.005805f
C32 cap_bsw_1/VPBT3 VDDA 0.858856f
C33 ncell_bsw_sw_1/VBOOT VSSA 0.040611f
C34 cap_bsw_1/VPBT2 VI 0.044479f
C35 cap_bsw_1/VPBT3 cap_bsw_1/VPBT2 0.037813f
C36 VI cap_bsw_1/VNBT3 -0.030413f
C37 cap_bsw_1/VPBT3 cap_bsw_1/VNBT3 0.45526f
C38 CLKS VI 0.059318f
C39 cap_bsw_1/VPBT3 CLKS 0.027275f
C40 VO ncell_bsw_sw_1/SWITCHING 0.038301f
C41 cap_bsw_1/VPBT3 ncell_bsw_dischrg_1/a_179_n1156# 0.015245f
C42 cap_bsw_1/VPBT1 ncell_bsw_sw_1/VBOOT 0.001455f
C43 CLKSB ncell_bsw_sw_1/SWITCHING 0.750737f
C44 cap_bsw_1/VPBT1 VSSA 0.181721f
C45 VDDA VO 4e-19
C46 cap_bsw_1/VPBT2 VO 0.039895f
C47 VDDA CLKSB 0.010193f
C48 VO cap_bsw_1/VNBT3 0.115938f
C49 CLKS VO 0.049474f
C50 CLKSB cap_bsw_1/VPBT2 0.977878f
C51 CLKSB cap_bsw_1/VNBT3 0.559164f
C52 CLKS CLKSB 1.268383f
C53 CLKSB ncell_bsw_dischrg_1/a_179_n1156# 1.21e-19
C54 cap_bsw_1/VPBT3 VI 0.008913f
C55 ncell_bsw_sw_1/VBOOT ncell_bsw_sw_1/SWITCHING 0.099269f
C56 VO VI 0.387392f
C57 cap_bsw_1/VPBT3 VO 0.003418f
C58 CLKSB VI 0.13119f
C59 cap_bsw_1/VPBT3 CLKSB 0.366048f
C60 VSSA ncell_bsw_sw_1/SWITCHING 0.08219f
C61 ncell_bsw_sw_1/VBOOT VDDA 0.589142f
C62 ncell_bsw_sw_1/VBOOT cap_bsw_1/VPBT2 0.002425f
C63 ncell_bsw_sw_1/VBOOT cap_bsw_1/VNBT3 0.379112f
C64 cap_bsw_1/VPBT1 ncell_bsw_sw_1/SWITCHING 0.511487f
C65 ncell_bsw_sw_1/VBOOT CLKS 0.017424f
C66 VDDA VSSA 0.41813f
C67 ncell_bsw_sw_1/VBOOT ncell_bsw_dischrg_1/a_179_n1156# 6.06e-21
C68 VSSA cap_bsw_1/VPBT2 0.065658f
C69 VSSA cap_bsw_1/VNBT3 0.109088f
C70 CLKS VSSA 0.063239f
C71 cap_bsw_1/VPBT1 VDDA 0.571642f
C72 CLKSB VO 0.070318f
C73 cap_bsw_1/VPBT1 0 1.693533f
C74 VDDA 0 1.933395f
C75 cap_bsw_1/VPBT2 0 1.444817f
C76 VSSA 0 -2.156982f
C77 ncell_bsw_dischrg_1/a_179_n1156# 0 0.072735f
C78 CLKSB 0 2.454724f
C79 cap_bsw_1/VNBT3 0 2.167416f
C80 VI 0 0.543435f
C81 ncell_bsw_sw_1/SWITCHING 0 1.559016f
C82 VO 0 0.101302f
C83 CLKS 0 1.132881f
C84 ncell_bsw_sw_1/VBOOT 0 2.030951f
C85 cap_bsw_1/VPBT3 0 2.856451f
.ends

