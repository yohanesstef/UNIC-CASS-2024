* NGSPICE file created from sh_bsw4.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_2XU92K a_n73_n100# w_n109_n162# a_15_n100# a_n15_n126#
+ VSUBS
X0 a_15_n100# a_n15_n126# a_n73_n100# w_n109_n162# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 w_n109_n162# a_15_n100# 0.006973f
C1 a_n15_n126# w_n109_n162# 0.022339f
C2 w_n109_n162# a_n73_n100# 0.006973f
C3 a_n15_n126# a_15_n100# 0.005542f
C4 a_15_n100# a_n73_n100# 0.162113f
C5 a_n15_n126# a_n73_n100# 0.005542f
C6 a_15_n100# VSUBS 0.111398f
C7 a_n73_n100# VSUBS 0.111398f
C8 a_n15_n126# VSUBS 0.043702f
C9 w_n109_n162# VSUBS 0.211896f
.ends

.subckt sky130_fd_pr__nfet_01v8_RH3MT7 a_n15_n76# a_n73_n50# a_15_n50# VSUBS
X0 a_15_n50# a_n15_n76# a_n73_n50# VSUBS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
C0 a_n73_n50# a_n15_n76# 0.003563f
C1 a_n15_n76# a_15_n50# 0.003563f
C2 a_n73_n50# a_15_n50# 0.082646f
C3 a_15_n50# VSUBS 0.076084f
C4 a_n73_n50# VSUBS 0.076084f
C5 a_n15_n76# VSUBS 0.066041f
.ends

.subckt inv_bsw IN OUT VPWR VPB VGND VNB
Xsky130_fd_pr__pfet_01v8_2XU92K_1 VPWR VPB OUT IN VNB sky130_fd_pr__pfet_01v8_2XU92K
Xsky130_fd_pr__nfet_01v8_RH3MT7_1 IN VGND OUT VNB sky130_fd_pr__nfet_01v8_RH3MT7
C0 VGND OUT 2.13e-19
C1 VGND IN 0.039434f
C2 VPB OUT 0.018962f
C3 IN VPB 0.032522f
C4 VPB VPWR 0.014235f
C5 IN OUT 0.037615f
C6 OUT VPWR 2.13e-19
C7 IN VPWR 0.040691f
C8 VGND VPB 1.03e-19
C9 VGND VNB 0.068517f
C10 OUT VNB 0.200334f
C11 VPWR VNB 0.090398f
C12 IN VNB 0.186801f
C13 VPB VNB 0.302938f
.ends

.subckt sky130_fd_pr__pfet_01v8_275TTJ a_n15_n76# w_n109_n112# a_n73_n50# a_15_n50#
+ VSUBS
X0 a_15_n50# a_n15_n76# a_n73_n50# w_n109_n112# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
C0 w_n109_n112# a_n73_n50# 0.00578f
C1 a_15_n50# a_n15_n76# 0.003563f
C2 w_n109_n112# a_15_n50# 0.00578f
C3 a_15_n50# a_n73_n50# 0.082646f
C4 w_n109_n112# a_n15_n76# 0.022339f
C5 a_n15_n76# a_n73_n50# 0.003563f
C6 a_15_n50# VSUBS 0.070304f
C7 a_n73_n50# VSUBS 0.070304f
C8 a_n15_n76# VSUBS 0.043702f
C9 w_n109_n112# VSUBS 0.146496f
.ends

.subckt pcell_bsw_dischrg VPBT3 SWITCHING VBOOT VSUBS
Xsky130_fd_pr__pfet_01v8_275TTJ_6 VPBT3 VPBT3 VPBT3 VBOOT VSUBS sky130_fd_pr__pfet_01v8_275TTJ
Xsky130_fd_pr__pfet_01v8_275TTJ_7 SWITCHING VPBT3 VPBT3 VBOOT VSUBS sky130_fd_pr__pfet_01v8_275TTJ
Xsky130_fd_pr__pfet_01v8_275TTJ_8 VPBT3 VPBT3 VBOOT VPBT3 VSUBS sky130_fd_pr__pfet_01v8_275TTJ
Xsky130_fd_pr__pfet_01v8_275TTJ_0 SWITCHING VPBT3 VBOOT VPBT3 VSUBS sky130_fd_pr__pfet_01v8_275TTJ
Xsky130_fd_pr__pfet_01v8_275TTJ_1 SWITCHING VPBT3 VPBT3 VBOOT VSUBS sky130_fd_pr__pfet_01v8_275TTJ
Xsky130_fd_pr__pfet_01v8_275TTJ_2 SWITCHING VPBT3 VBOOT VPBT3 VSUBS sky130_fd_pr__pfet_01v8_275TTJ
Xsky130_fd_pr__pfet_01v8_275TTJ_3 VPBT3 VPBT3 VPBT3 VBOOT VSUBS sky130_fd_pr__pfet_01v8_275TTJ
Xsky130_fd_pr__pfet_01v8_275TTJ_4 VPBT3 VPBT3 VBOOT VPBT3 VSUBS sky130_fd_pr__pfet_01v8_275TTJ
C0 VPBT3 SWITCHING 0.305567f
C1 VBOOT SWITCHING 0.044932f
C2 VPBT3 VBOOT 0.175809f
C3 VBOOT VSUBS 0.230584f
C4 VPBT3 VSUBS 1.939276f
C5 SWITCHING VSUBS 0.110218f
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_UCPR8Z m3_n386_n240# c1_n346_n200# VSUBS
X0 c1_n346_n200# m3_n386_n240# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
C0 c1_n346_n200# m3_n386_n240# 0.507132f
C1 c1_n346_n200# VSUBS 0.169673f
C2 m3_n386_n240# VSUBS 0.762748f
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_VCTT89 m3_n386_n240# c1_n346_n200# VSUBS
X0 c1_n346_n200# m3_n386_n240# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
C0 c1_n346_n200# m3_n386_n240# 0.507132f
C1 c1_n346_n200# VSUBS 0.169673f
C2 m3_n386_n240# VSUBS 0.762748f
.ends

.subckt cap_bsw VPBT1 VNBT1 VPBT2 VPBT3 VNBT3 CLKS VSUBS
Xsky130_fd_pr__cap_mim_m3_1_UCPR8Z_0 VNBT1 VPBT1 VSUBS sky130_fd_pr__cap_mim_m3_1_UCPR8Z
Xsky130_fd_pr__cap_mim_m3_1_VCTT89_0 VNBT3 VPBT3 VSUBS sky130_fd_pr__cap_mim_m3_1_VCTT89
Xsky130_fd_pr__cap_mim_m3_1_VCTT89_1 VNBT3 VPBT3 VSUBS sky130_fd_pr__cap_mim_m3_1_VCTT89
XXC2 CLKS VPBT2 VSUBS sky130_fd_pr__cap_mim_m3_1_VCTT89
C0 VNBT3 CLKS 0.312674f
C1 CLKS VPBT3 0.13591f
C2 CLKS VNBT1 0.382401f
C3 CLKS VPBT1 0.012183f
C4 VNBT3 VPBT3 0.143473f
C5 VNBT3 VNBT1 0.312674f
C6 VPBT2 VNBT1 0.012183f
C7 VNBT1 VPBT3 0.13591f
C8 VPBT2 VPBT1 0.084078f
C9 VPBT3 VSUBS 0.160558f
C10 VNBT3 VSUBS 1.011946f
C11 VPBT2 VSUBS 0.11587f
C12 CLKS VSUBS 0.424282f
C13 VPBT1 VSUBS 0.11587f
C14 VNBT1 VSUBS 0.424282f
.ends

.subckt sky130_fd_pr__nfet_01v8_QS6TK8 a_30_n50# a_n30_n76# a_n88_n50# VSUBS
X0 a_30_n50# a_n30_n76# a_n88_n50# VSUBS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.3
C0 a_n88_n50# a_30_n50# 0.061754f
C1 a_n30_n76# a_n88_n50# 0.006618f
C2 a_n30_n76# a_30_n50# 0.006618f
C3 a_30_n50# VSUBS 0.076817f
C4 a_n88_n50# VSUBS 0.076817f
C5 a_n30_n76# VSUBS 0.103343f
.ends

.subckt sky130_fd_pr__nfet_01v8_6J3TAM a_n15_n76# a_n73_n50# a_15_n50# VSUBS
X0 a_15_n50# a_n15_n76# a_n73_n50# VSUBS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
C0 a_n73_n50# a_15_n50# 0.082646f
C1 a_n15_n76# a_n73_n50# 0.003563f
C2 a_n15_n76# a_15_n50# 0.003563f
C3 a_15_n50# VSUBS 0.076084f
C4 a_n73_n50# VSUBS 0.076084f
C5 a_n15_n76# VSUBS 0.066041f
.ends

.subckt ncell_bsw_sw VI VBOOT VNBT1 VNBT3 SWITCHING VSSA VO
Xsky130_fd_pr__nfet_01v8_QS6TK8_0 VI VBOOT VNBT3 VSSA sky130_fd_pr__nfet_01v8_QS6TK8
Xsky130_fd_pr__nfet_01v8_QS6TK8_1 VO VBOOT VI VSSA sky130_fd_pr__nfet_01v8_QS6TK8
Xsky130_fd_pr__nfet_01v8_QS6TK8_2 VI VBOOT VO VSSA sky130_fd_pr__nfet_01v8_QS6TK8
Xsky130_fd_pr__nfet_01v8_QS6TK8_4 VI VI VI VSSA sky130_fd_pr__nfet_01v8_QS6TK8
Xsky130_fd_pr__nfet_01v8_QS6TK8_3 VNBT3 VBOOT VI VSSA sky130_fd_pr__nfet_01v8_QS6TK8
Xsky130_fd_pr__nfet_01v8_6J3TAM_10 SWITCHING SWITCHING SWITCHING VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_QS6TK8_5 VI VI VI VSSA sky130_fd_pr__nfet_01v8_QS6TK8
Xsky130_fd_pr__nfet_01v8_QS6TK8_6 VO VBOOT VI VSSA sky130_fd_pr__nfet_01v8_QS6TK8
Xsky130_fd_pr__nfet_01v8_QS6TK8_7 VI VBOOT VO VSSA sky130_fd_pr__nfet_01v8_QS6TK8
Xsky130_fd_pr__nfet_01v8_6J3TAM_0 VBOOT SWITCHING VNBT3 VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_1 VBOOT VNBT3 SWITCHING VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_2 VNBT1 VSSA VNBT3 VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_3 VNBT1 VNBT3 VSSA VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_4 VSSA VSSA VSSA VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_5 VSSA VSSA VSSA VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_6 SWITCHING SWITCHING SWITCHING VSSA sky130_fd_pr__nfet_01v8_6J3TAM
C0 VI VSSA 0.003263f
C1 VO VSSA -3.54e-19
C2 VBOOT VNBT3 0.312731f
C3 VI SWITCHING 0.007828f
C4 VO SWITCHING 2.07e-19
C5 VNBT1 VSSA 0.161521f
C6 VBOOT VI 0.383013f
C7 VNBT1 SWITCHING 0.08682f
C8 VBOOT VO 0.051806f
C9 VI VNBT3 0.543276f
C10 VO VNBT3 0.032599f
C11 VBOOT VNBT1 0.116444f
C12 VNBT1 VNBT3 0.39543f
C13 VI VO 0.292146f
C14 SWITCHING VSSA 0.147075f
C15 VI VNBT1 0.189617f
C16 VBOOT VSSA -0.009935f
C17 VNBT1 VO 0.028509f
C18 VBOOT SWITCHING 0.135406f
C19 VSSA VNBT3 0.021985f
C20 SWITCHING VNBT3 0.007802f
C21 VNBT3 0 0.430447f
C22 VSSA 0 0.357545f
C23 VNBT1 0 0.663646f
C24 SWITCHING 0 0.56538f
C25 VO 0 0.044245f
C26 VBOOT 0 0.941026f
C27 VI 0 0.676943f
.ends

.subckt ncell_bsw_dischrg VDDA CLKSB VBOOT VSSA a_179_n1156#
Xsky130_fd_pr__nfet_01v8_6J3TAM_0 VBOOT VBOOT VBOOT VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_1 VSSA VSSA VSSA VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_2 CLKSB VSSA a_179_n1156# VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_3 VDDA a_179_n1156# VBOOT VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_4 VBOOT VBOOT VBOOT VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_5 VDDA VBOOT a_179_n1156# VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_6 CLKSB a_179_n1156# VSSA VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_7 VSSA VSSA VSSA VSSA sky130_fd_pr__nfet_01v8_6J3TAM
C0 VDDA VSSA 0.022289f
C1 a_179_n1156# VSSA -0.001926f
C2 VBOOT CLKSB 0.336066f
C3 VDDA VBOOT 0.108129f
C4 a_179_n1156# VBOOT 0.003556f
C5 VBOOT VSSA 0.132444f
C6 VDDA CLKSB 0.09168f
C7 a_179_n1156# CLKSB 0.135282f
C8 CLKSB VSSA 0.049316f
C9 a_179_n1156# VDDA 0.08975f
C10 VSSA 0 0.030694f
C11 a_179_n1156# 0 0.084125f
C12 CLKSB 0 0.561057f
C13 VBOOT 0 1.039818f
C14 VDDA 0 0.348624f
.ends

.subckt ncell_bsw VDDA VPBT1 VPBT2 VPBT3 VSSA
Xsky130_fd_pr__nfet_01v8_6J3TAM_10 VPBT1 VDDA VPBT3 VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_11 VPBT1 VPBT1 VPBT1 VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_12 VPBT2 VDDA VPBT1 VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_13 VPBT1 VPBT2 VDDA VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_14 VPBT2 VPBT2 VPBT2 VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_15 VPBT1 VPBT1 VPBT1 VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_0 VDDA VDDA VDDA VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_1 VPBT1 VPBT2 VDDA VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_2 VPBT2 VDDA VPBT1 VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_3 VPBT2 VPBT2 VPBT2 VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_4 VPBT3 VPBT3 VPBT3 VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_5 VPBT1 VPBT3 VDDA VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_6 VDDA VDDA VDDA VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_7 VPBT3 VPBT3 VPBT3 VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_8 VDDA VDDA VDDA VSSA sky130_fd_pr__nfet_01v8_6J3TAM
Xsky130_fd_pr__nfet_01v8_6J3TAM_9 VDDA VDDA VDDA VSSA sky130_fd_pr__nfet_01v8_6J3TAM
C0 VPBT2 VDDA 0.291541f
C1 VPBT2 VPBT1 0.461288f
C2 VPBT1 VDDA 0.670526f
C3 VPBT3 VPBT2 0.238169f
C4 VPBT3 VDDA 0.357952f
C5 VPBT3 VPBT1 0.427097f
C6 VDDA VSSA 0.682311f
C7 VPBT3 VSSA 0.54034f
C8 VPBT1 VSSA 1.406676f
C9 VPBT2 VSSA 1.405102f
.ends

.subckt sh_bsw3 ncell_bsw_dischrg_0/VDDA ncell_bsw_dischrg_0/a_179_n1156# inv_bsw_0/OUT
+ inv_bsw_0/IN inv_bsw_0/VPB ncell_bsw_sw_1/VO ncell_bsw_sw_1/VI cap_bsw_1/VPBT3 cap_bsw_1/VPBT2
+ inv_bsw_0/VGND cap_bsw_1/VNBT1 cap_bsw_1/VPBT1 inv_bsw_0/VPWR ncell_bsw_sw_1/VBOOT
+ VSUBS
Xinv_bsw_0 inv_bsw_0/IN inv_bsw_0/OUT inv_bsw_0/VPWR inv_bsw_0/VPB inv_bsw_0/VGND
+ VSUBS inv_bsw
Xpcell_bsw_dischrg_0 cap_bsw_1/VPBT3 inv_bsw_0/OUT ncell_bsw_sw_1/VBOOT VSUBS pcell_bsw_dischrg
Xcap_bsw_1 cap_bsw_1/VPBT1 cap_bsw_1/VNBT1 cap_bsw_1/VPBT2 cap_bsw_1/VPBT3 inv_bsw_0/VGND
+ inv_bsw_0/IN VSUBS cap_bsw
Xncell_bsw_sw_1 ncell_bsw_sw_1/VI ncell_bsw_sw_1/VBOOT cap_bsw_1/VNBT1 inv_bsw_0/VGND
+ inv_bsw_0/OUT VSUBS ncell_bsw_sw_1/VO ncell_bsw_sw
Xncell_bsw_dischrg_0 ncell_bsw_dischrg_0/VDDA cap_bsw_1/VNBT1 ncell_bsw_sw_1/VBOOT
+ VSUBS ncell_bsw_dischrg_0/a_179_n1156# ncell_bsw_dischrg
Xncell_bsw_1 inv_bsw_0/VPWR cap_bsw_1/VPBT1 cap_bsw_1/VPBT2 cap_bsw_1/VPBT3 VSUBS
+ ncell_bsw
C0 inv_bsw_0/OUT cap_bsw_1/VPBT1 0.043726f
C1 inv_bsw_0/VPB ncell_bsw_sw_1/VI 4.15e-21
C2 ncell_bsw_sw_1/VI cap_bsw_1/VPBT3 0.001756f
C3 cap_bsw_1/VNBT1 ncell_bsw_dischrg_0/VDDA 9.38e-19
C4 ncell_bsw_dischrg_0/a_179_n1156# ncell_bsw_sw_1/VI 1.8e-20
C5 ncell_bsw_sw_1/VO ncell_bsw_dischrg_0/VDDA 4.97e-20
C6 inv_bsw_0/VPWR inv_bsw_0/IN 0.169569f
C7 inv_bsw_0/VGND inv_bsw_0/IN 6.12e-19
C8 inv_bsw_0/OUT cap_bsw_1/VNBT1 0.680974f
C9 inv_bsw_0/OUT ncell_bsw_sw_1/VO 0.034792f
C10 inv_bsw_0/VPB VSUBS 0.013335f
C11 VSUBS cap_bsw_1/VPBT3 0.295196f
C12 ncell_bsw_dischrg_0/a_179_n1156# VSUBS 0.005616f
C13 inv_bsw_0/VPWR cap_bsw_1/VPBT2 0.229682f
C14 inv_bsw_0/VGND cap_bsw_1/VPBT2 0.903526f
C15 inv_bsw_0/VPB cap_bsw_1/VPBT3 8.49e-20
C16 ncell_bsw_sw_1/VBOOT inv_bsw_0/VPWR 0.003532f
C17 inv_bsw_0/VGND ncell_bsw_sw_1/VBOOT 0.35759f
C18 inv_bsw_0/OUT inv_bsw_0/IN 0.019226f
C19 ncell_bsw_sw_1/VI inv_bsw_0/VPWR 1.89e-20
C20 ncell_bsw_sw_1/VI inv_bsw_0/VGND 0.120248f
C21 ncell_bsw_sw_1/VBOOT ncell_bsw_dischrg_0/VDDA 0.001697f
C22 inv_bsw_0/OUT cap_bsw_1/VPBT2 0.067211f
C23 VSUBS inv_bsw_0/VPWR 0.011986f
C24 inv_bsw_0/OUT ncell_bsw_sw_1/VBOOT 0.188704f
C25 VSUBS inv_bsw_0/VGND 0.307046f
C26 cap_bsw_1/VNBT1 cap_bsw_1/VPBT1 0.314337f
C27 ncell_bsw_sw_1/VI ncell_bsw_dischrg_0/VDDA 3.28e-19
C28 ncell_bsw_sw_1/VO cap_bsw_1/VPBT1 1.11e-20
C29 inv_bsw_0/VPB inv_bsw_0/VPWR 0.009513f
C30 inv_bsw_0/VPWR cap_bsw_1/VPBT3 0.025386f
C31 inv_bsw_0/VPB inv_bsw_0/VGND 4.69e-19
C32 ncell_bsw_sw_1/VI inv_bsw_0/OUT 0.270848f
C33 inv_bsw_0/VGND cap_bsw_1/VPBT3 0.41275f
C34 ncell_bsw_dischrg_0/a_179_n1156# inv_bsw_0/VGND 1.57e-20
C35 ncell_bsw_sw_1/VO cap_bsw_1/VNBT1 0.018792f
C36 VSUBS ncell_bsw_dischrg_0/VDDA 0.002527f
C37 inv_bsw_0/IN cap_bsw_1/VPBT1 0.155073f
C38 VSUBS inv_bsw_0/OUT 0.19398f
C39 inv_bsw_0/VPB inv_bsw_0/OUT 3.23e-20
C40 inv_bsw_0/IN cap_bsw_1/VNBT1 0.324472f
C41 inv_bsw_0/OUT cap_bsw_1/VPBT3 0.360643f
C42 ncell_bsw_dischrg_0/a_179_n1156# inv_bsw_0/OUT 0.003454f
C43 ncell_bsw_sw_1/VO inv_bsw_0/IN 2.66e-19
C44 cap_bsw_1/VPBT2 cap_bsw_1/VPBT1 0.321807f
C45 ncell_bsw_sw_1/VBOOT cap_bsw_1/VPBT1 0.00177f
C46 inv_bsw_0/VGND inv_bsw_0/VPWR 0.068416f
C47 cap_bsw_1/VNBT1 cap_bsw_1/VPBT2 0.018862f
C48 ncell_bsw_sw_1/VI cap_bsw_1/VPBT1 1.74e-19
C49 ncell_bsw_sw_1/VO cap_bsw_1/VPBT2 3.54e-19
C50 ncell_bsw_sw_1/VBOOT cap_bsw_1/VNBT1 0.578002f
C51 ncell_bsw_sw_1/VBOOT ncell_bsw_sw_1/VO 0.006678f
C52 inv_bsw_0/VGND ncell_bsw_dischrg_0/VDDA 2.75e-19
C53 ncell_bsw_sw_1/VI cap_bsw_1/VNBT1 0.11536f
C54 VSUBS cap_bsw_1/VPBT1 0.017379f
C55 ncell_bsw_sw_1/VI ncell_bsw_sw_1/VO 0.357567f
C56 inv_bsw_0/OUT inv_bsw_0/VPWR 0.06661f
C57 inv_bsw_0/OUT inv_bsw_0/VGND 1.377584f
C58 inv_bsw_0/IN cap_bsw_1/VPBT2 0.225363f
C59 inv_bsw_0/VPB cap_bsw_1/VPBT1 0.009776f
C60 ncell_bsw_sw_1/VBOOT inv_bsw_0/IN 0.004329f
C61 cap_bsw_1/VPBT1 cap_bsw_1/VPBT3 0.220569f
C62 VSUBS cap_bsw_1/VNBT1 0.048945f
C63 VSUBS ncell_bsw_sw_1/VO 5.04e-19
C64 ncell_bsw_sw_1/VI inv_bsw_0/IN 0.002078f
C65 inv_bsw_0/OUT ncell_bsw_dischrg_0/VDDA 0.001209f
C66 inv_bsw_0/VPB cap_bsw_1/VNBT1 0.001291f
C67 cap_bsw_1/VNBT1 cap_bsw_1/VPBT3 0.120821f
C68 ncell_bsw_sw_1/VBOOT cap_bsw_1/VPBT2 0.002328f
C69 ncell_bsw_sw_1/VO cap_bsw_1/VPBT3 2.84e-20
C70 ncell_bsw_dischrg_0/a_179_n1156# cap_bsw_1/VNBT1 1.45e-19
C71 ncell_bsw_dischrg_0/a_179_n1156# ncell_bsw_sw_1/VO 8.69e-21
C72 VSUBS inv_bsw_0/IN 0.02742f
C73 ncell_bsw_sw_1/VI cap_bsw_1/VPBT2 0.002409f
C74 ncell_bsw_sw_1/VI ncell_bsw_sw_1/VBOOT 0.308781f
C75 inv_bsw_0/VPB inv_bsw_0/IN 0.027914f
C76 inv_bsw_0/IN cap_bsw_1/VPBT3 0.045769f
C77 inv_bsw_0/VPWR cap_bsw_1/VPBT1 0.029276f
C78 inv_bsw_0/VGND cap_bsw_1/VPBT1 0.134697f
C79 VSUBS cap_bsw_1/VPBT2 0.025899f
C80 VSUBS ncell_bsw_sw_1/VBOOT 0.261316f
C81 inv_bsw_0/VPWR cap_bsw_1/VNBT1 0.005906f
C82 inv_bsw_0/VGND cap_bsw_1/VNBT1 0.236762f
C83 inv_bsw_0/VPB cap_bsw_1/VPBT2 0.008099f
C84 cap_bsw_1/VPBT2 cap_bsw_1/VPBT3 0.144957f
C85 inv_bsw_0/VGND ncell_bsw_sw_1/VO 0.055948f
C86 ncell_bsw_sw_1/VI VSUBS 0.003132f
C87 ncell_bsw_sw_1/VBOOT cap_bsw_1/VPBT3 0.689421f
C88 ncell_bsw_dischrg_0/a_179_n1156# ncell_bsw_sw_1/VBOOT 8.09e-19
C89 inv_bsw_0/VPWR 0 0.733294f
C90 cap_bsw_1/VPBT3 0 2.519834f
C91 cap_bsw_1/VPBT1 0 2.045305f
C92 cap_bsw_1/VPBT2 0 1.332593f
C93 ncell_bsw_dischrg_0/a_179_n1156# 0 0.084125f
C94 ncell_bsw_dischrg_0/VDDA 0 0.348624f
C95 inv_bsw_0/VGND 0 1.846506f
C96 VSUBS 0 -1.57265f
C97 cap_bsw_1/VNBT1 0 2.833024f
C98 inv_bsw_0/OUT 0 0.977822f
C99 ncell_bsw_sw_1/VO 0 0.070107f
C100 ncell_bsw_sw_1/VI 0 0.756526f
C101 ncell_bsw_sw_1/VBOOT 0 2.465944f
C102 inv_bsw_0/IN 0 0.650316f
C103 inv_bsw_0/VPB 0 0.304109f
.ends

.subckt sh_bsw4 VDDA CLKS CLKSB VIP VIN VSSA VCP VCN
Xsh_bsw3_0 VDDA sh_bsw3_0/ncell_bsw_dischrg_0/a_179_n1156# sh_bsw3_0/inv_bsw_0/OUT
+ CLKS VDDA VCP VIP sh_bsw3_0/cap_bsw_1/VPBT3 sh_bsw3_0/cap_bsw_1/VPBT2 sh_bsw3_0/inv_bsw_0/VGND
+ CLKSB sh_bsw3_0/cap_bsw_1/VPBT1 VDDA sh_bsw3_0/ncell_bsw_sw_1/VBOOT VSSA sh_bsw3
Xsh_bsw3_1 VDDA sh_bsw3_1/ncell_bsw_dischrg_0/a_179_n1156# sh_bsw3_1/inv_bsw_0/OUT
+ CLKS VDDA VCN VIN sh_bsw3_1/cap_bsw_1/VPBT3 sh_bsw3_1/cap_bsw_1/VPBT2 sh_bsw3_1/inv_bsw_0/VGND
+ CLKSB sh_bsw3_1/cap_bsw_1/VPBT1 VDDA sh_bsw3_1/ncell_bsw_sw_1/VBOOT VSSA sh_bsw3
C0 VIN sh_bsw3_0/ncell_bsw_sw_1/VBOOT 0.001272f
C1 sh_bsw3_1/ncell_bsw_sw_1/VBOOT CLKSB -0.107908f
C2 VSSA sh_bsw3_0/inv_bsw_0/OUT 0.005537f
C3 sh_bsw3_0/inv_bsw_0/VGND CLKS 0.457889f
C4 sh_bsw3_0/ncell_bsw_dischrg_0/a_179_n1156# sh_bsw3_1/cap_bsw_1/VPBT1 2.37e-20
C5 sh_bsw3_1/ncell_bsw_dischrg_0/a_179_n1156# VDDA 0.026945f
C6 VCP VCN 0.002064f
C7 sh_bsw3_1/cap_bsw_1/VPBT2 CLKS -0.003521f
C8 CLKSB VDDA 2.752979f
C9 sh_bsw3_1/ncell_bsw_dischrg_0/a_179_n1156# sh_bsw3_1/inv_bsw_0/VGND -3.3e-21
C10 CLKSB VIP -0.00374f
C11 CLKS sh_bsw3_1/cap_bsw_1/VPBT1 -0.010271f
C12 CLKSB sh_bsw3_1/inv_bsw_0/VGND 0.387797f
C13 CLKS sh_bsw3_0/cap_bsw_1/VPBT1 0.14811f
C14 CLKSB sh_bsw3_1/cap_bsw_1/VPBT3 0.051241f
C15 CLKS VCN 0.036131f
C16 CLKSB sh_bsw3_0/cap_bsw_1/VPBT3 0.004275f
C17 sh_bsw3_1/ncell_bsw_sw_1/VBOOT sh_bsw3_0/inv_bsw_0/OUT 0.023472f
C18 VIN VCN -0.002452f
C19 sh_bsw3_0/cap_bsw_1/VPBT2 VSSA 9.83e-19
C20 VDDA sh_bsw3_0/inv_bsw_0/OUT 0.038729f
C21 VIN CLKS 0.153993f
C22 sh_bsw3_1/ncell_bsw_sw_1/VBOOT VSSA 0.028502f
C23 sh_bsw3_1/inv_bsw_0/VGND sh_bsw3_0/inv_bsw_0/OUT 5.9e-21
C24 sh_bsw3_1/inv_bsw_0/OUT CLKSB -0.185069f
C25 VDDA VSSA 0.197733f
C26 sh_bsw3_1/cap_bsw_1/VPBT3 sh_bsw3_0/inv_bsw_0/OUT 0.002417f
C27 VIP VSSA 2.22e-20
C28 VSSA sh_bsw3_1/inv_bsw_0/VGND 0.078768f
C29 CLKSB sh_bsw3_0/ncell_bsw_sw_1/VBOOT -0.151631f
C30 sh_bsw3_1/ncell_bsw_sw_1/VBOOT sh_bsw3_0/cap_bsw_1/VPBT2 0.017562f
C31 VSSA sh_bsw3_1/cap_bsw_1/VPBT3 0.074997f
C32 sh_bsw3_0/inv_bsw_0/VGND CLKSB 0.002724f
C33 sh_bsw3_1/cap_bsw_1/VPBT2 CLKSB 0.038006f
C34 sh_bsw3_0/cap_bsw_1/VPBT2 VDDA 0.08244f
C35 VSSA sh_bsw3_0/cap_bsw_1/VPBT3 0.08109f
C36 VCP CLKSB -0.00315f
C37 sh_bsw3_1/ncell_bsw_dischrg_0/a_179_n1156# sh_bsw3_0/cap_bsw_1/VPBT1 2.37e-20
C38 sh_bsw3_1/inv_bsw_0/OUT sh_bsw3_0/inv_bsw_0/OUT 0.004582f
C39 sh_bsw3_1/ncell_bsw_sw_1/VBOOT VDDA 0.218522f
C40 CLKSB sh_bsw3_1/cap_bsw_1/VPBT1 0.131505f
C41 CLKSB sh_bsw3_0/cap_bsw_1/VPBT1 -0.024801f
C42 sh_bsw3_1/ncell_bsw_sw_1/VBOOT VIP 0.001272f
C43 sh_bsw3_1/ncell_bsw_sw_1/VBOOT sh_bsw3_1/inv_bsw_0/VGND -4.62e-19
C44 sh_bsw3_0/cap_bsw_1/VPBT2 sh_bsw3_1/cap_bsw_1/VPBT3 5.19e-21
C45 sh_bsw3_1/ncell_bsw_dischrg_0/a_179_n1156# VCN -1.83e-21
C46 sh_bsw3_0/ncell_bsw_dischrg_0/a_179_n1156# CLKSB 1.29e-19
C47 sh_bsw3_0/cap_bsw_1/VPBT2 sh_bsw3_0/cap_bsw_1/VPBT3 -5.69e-20
C48 CLKSB VCN -0.006138f
C49 sh_bsw3_1/inv_bsw_0/OUT VSSA 0.082687f
C50 VDDA VIP 0.00751f
C51 sh_bsw3_1/ncell_bsw_sw_1/VBOOT sh_bsw3_1/cap_bsw_1/VPBT3 6.25e-31
C52 VDDA sh_bsw3_1/inv_bsw_0/VGND 0.144446f
C53 CLKS sh_bsw3_1/ncell_bsw_dischrg_0/a_179_n1156# 1.81e-19
C54 sh_bsw3_1/ncell_bsw_sw_1/VBOOT sh_bsw3_0/cap_bsw_1/VPBT3 0.098391f
C55 VIN sh_bsw3_1/ncell_bsw_dischrg_0/a_179_n1156# -3.78e-21
C56 CLKSB CLKS 1.794579f
C57 VDDA sh_bsw3_1/cap_bsw_1/VPBT3 0.003333f
C58 sh_bsw3_0/ncell_bsw_sw_1/VBOOT VSSA -0.00746f
C59 VIN CLKSB -0.071375f
C60 VDDA sh_bsw3_0/cap_bsw_1/VPBT3 0.003438f
C61 sh_bsw3_1/cap_bsw_1/VPBT1 sh_bsw3_0/inv_bsw_0/OUT 3.83e-20
C62 VIP sh_bsw3_1/cap_bsw_1/VPBT3 0.00545f
C63 sh_bsw3_1/inv_bsw_0/VGND sh_bsw3_1/cap_bsw_1/VPBT3 -3.07e-19
C64 sh_bsw3_0/cap_bsw_1/VPBT1 sh_bsw3_0/inv_bsw_0/OUT 3.55e-33
C65 sh_bsw3_0/inv_bsw_0/VGND VSSA 0.072739f
C66 sh_bsw3_1/cap_bsw_1/VPBT2 VSSA 0.003362f
C67 sh_bsw3_0/cap_bsw_1/VPBT3 sh_bsw3_1/inv_bsw_0/VGND 0.004489f
C68 sh_bsw3_1/ncell_bsw_sw_1/VBOOT sh_bsw3_1/inv_bsw_0/OUT -0.00263f
C69 sh_bsw3_0/cap_bsw_1/VPBT3 sh_bsw3_1/cap_bsw_1/VPBT3 0.071805f
C70 VSSA sh_bsw3_1/cap_bsw_1/VPBT1 0.006382f
C71 sh_bsw3_0/cap_bsw_1/VPBT1 VSSA 0.005715f
C72 sh_bsw3_1/inv_bsw_0/OUT VDDA 0.015728f
C73 CLKS sh_bsw3_0/inv_bsw_0/OUT 1.82e-21
C74 sh_bsw3_0/inv_bsw_0/VGND sh_bsw3_0/cap_bsw_1/VPBT2 -0.001907f
C75 sh_bsw3_1/ncell_bsw_sw_1/VBOOT sh_bsw3_0/ncell_bsw_sw_1/VBOOT 0.109577f
C76 VSSA VCN 0.008016f
C77 sh_bsw3_0/inv_bsw_0/VGND sh_bsw3_1/ncell_bsw_sw_1/VBOOT 0.290604f
C78 sh_bsw3_0/ncell_bsw_sw_1/VBOOT VDDA 0.374667f
C79 CLKS VSSA 0.260693f
C80 sh_bsw3_0/cap_bsw_1/VPBT2 sh_bsw3_0/cap_bsw_1/VPBT1 -0.00753f
C81 sh_bsw3_0/ncell_bsw_sw_1/VBOOT VIP -5.68e-32
C82 VCP sh_bsw3_1/ncell_bsw_sw_1/VBOOT 8.12e-20
C83 sh_bsw3_0/inv_bsw_0/VGND VDDA 0.15279f
C84 sh_bsw3_0/ncell_bsw_sw_1/VBOOT sh_bsw3_1/inv_bsw_0/VGND 0.290602f
C85 sh_bsw3_1/inv_bsw_0/OUT sh_bsw3_0/cap_bsw_1/VPBT3 0.002417f
C86 VIN VSSA 0.010973f
C87 sh_bsw3_1/cap_bsw_1/VPBT2 VDDA 0.080136f
C88 sh_bsw3_1/ncell_bsw_sw_1/VBOOT sh_bsw3_0/cap_bsw_1/VPBT1 5.36e-19
C89 sh_bsw3_0/inv_bsw_0/VGND sh_bsw3_1/inv_bsw_0/VGND 0.006566f
C90 sh_bsw3_0/ncell_bsw_sw_1/VBOOT sh_bsw3_1/cap_bsw_1/VPBT3 0.098391f
C91 VCP VDDA 0.005992f
C92 sh_bsw3_1/cap_bsw_1/VPBT2 sh_bsw3_1/inv_bsw_0/VGND -0.001907f
C93 sh_bsw3_0/ncell_bsw_sw_1/VBOOT sh_bsw3_0/cap_bsw_1/VPBT3 1.14e-30
C94 VDDA sh_bsw3_1/cap_bsw_1/VPBT1 0.017836f
C95 CLKSB sh_bsw3_1/ncell_bsw_dischrg_0/a_179_n1156# -3.97e-20
C96 VDDA sh_bsw3_0/cap_bsw_1/VPBT1 0.018724f
C97 sh_bsw3_0/inv_bsw_0/VGND sh_bsw3_1/cap_bsw_1/VPBT3 0.004489f
C98 sh_bsw3_1/ncell_bsw_sw_1/VBOOT VCN -8.91e-21
C99 CLKS sh_bsw3_0/cap_bsw_1/VPBT2 0.035775f
C100 sh_bsw3_1/cap_bsw_1/VPBT2 sh_bsw3_1/cap_bsw_1/VPBT3 -5.66e-20
C101 sh_bsw3_0/inv_bsw_0/VGND sh_bsw3_0/cap_bsw_1/VPBT3 -3.07e-19
C102 sh_bsw3_0/ncell_bsw_dischrg_0/a_179_n1156# VDDA 0.031343f
C103 sh_bsw3_1/inv_bsw_0/VGND sh_bsw3_1/cap_bsw_1/VPBT1 -4.17e-19
C104 sh_bsw3_1/cap_bsw_1/VPBT2 sh_bsw3_0/cap_bsw_1/VPBT3 5.19e-21
C105 sh_bsw3_1/ncell_bsw_sw_1/VBOOT CLKS 0.03284f
C106 VDDA VCN 1.06e-20
C107 VIN sh_bsw3_1/ncell_bsw_sw_1/VBOOT -7.38e-20
C108 sh_bsw3_1/cap_bsw_1/VPBT1 sh_bsw3_1/cap_bsw_1/VPBT3 -9.04e-19
C109 sh_bsw3_0/cap_bsw_1/VPBT1 sh_bsw3_1/cap_bsw_1/VPBT3 0.001302f
C110 VCN sh_bsw3_1/inv_bsw_0/VGND -1.42e-32
C111 sh_bsw3_0/cap_bsw_1/VPBT3 sh_bsw3_1/cap_bsw_1/VPBT1 0.001302f
C112 CLKS VDDA 0.200137f
C113 sh_bsw3_1/inv_bsw_0/OUT sh_bsw3_0/ncell_bsw_sw_1/VBOOT 0.023472f
C114 sh_bsw3_0/cap_bsw_1/VPBT1 sh_bsw3_0/cap_bsw_1/VPBT3 -9.06e-19
C115 VIN VDDA 8.53e-20
C116 CLKS VIP -1.3e-21
C117 CLKS sh_bsw3_1/inv_bsw_0/VGND 0.179072f
C118 sh_bsw3_0/inv_bsw_0/VGND sh_bsw3_1/inv_bsw_0/OUT 5.9e-21
C119 VIN VIP 0.004361f
C120 CLKSB sh_bsw3_0/inv_bsw_0/OUT -0.01691f
C121 CLKS sh_bsw3_1/cap_bsw_1/VPBT3 1.17e-19
C122 CLKS sh_bsw3_0/cap_bsw_1/VPBT3 0.047194f
C123 sh_bsw3_1/cap_bsw_1/VPBT2 sh_bsw3_0/ncell_bsw_sw_1/VBOOT 0.017562f
C124 sh_bsw3_1/inv_bsw_0/OUT sh_bsw3_0/cap_bsw_1/VPBT1 3.83e-20
C125 VIN sh_bsw3_0/cap_bsw_1/VPBT3 0.00545f
C126 sh_bsw3_1/ncell_bsw_dischrg_0/a_179_n1156# VSSA -3.62e-19
C127 CLKSB VSSA 1.69037f
C128 sh_bsw3_0/ncell_bsw_sw_1/VBOOT sh_bsw3_1/cap_bsw_1/VPBT1 5.36e-19
C129 sh_bsw3_0/ncell_bsw_dischrg_0/a_179_n1156# sh_bsw3_0/ncell_bsw_sw_1/VBOOT -1.38e-19
C130 sh_bsw3_1/inv_bsw_0/OUT CLKS 0.270851f
C131 sh_bsw3_1/cap_bsw_1/VPBT2 sh_bsw3_1/cap_bsw_1/VPBT1 -0.00753f
C132 sh_bsw3_0/inv_bsw_0/VGND sh_bsw3_0/cap_bsw_1/VPBT1 -4.17e-19
C133 sh_bsw3_0/ncell_bsw_sw_1/VBOOT VCN 8.12e-20
C134 CLKSB sh_bsw3_0/cap_bsw_1/VPBT2 0.001253f
C135 sh_bsw3_1/ncell_bsw_sw_1/VBOOT sh_bsw3_1/ncell_bsw_dischrg_0/a_179_n1156# -3.1e-19
C136 CLKS sh_bsw3_0/ncell_bsw_sw_1/VBOOT 5.86e-20
C137 VDDA 0 4.053378f
C138 sh_bsw3_1/cap_bsw_1/VPBT3 0 2.519834f
C139 sh_bsw3_1/cap_bsw_1/VPBT1 0 2.045305f
C140 sh_bsw3_1/cap_bsw_1/VPBT2 0 1.332593f
C141 sh_bsw3_1/ncell_bsw_dischrg_0/a_179_n1156# 0 0.084125f
C142 sh_bsw3_1/inv_bsw_0/VGND 0 1.846506f
C143 VSSA 0 -2.423629f
C144 CLKSB 0 5.758368f
C145 sh_bsw3_1/inv_bsw_0/OUT 0 0.977822f
C146 VCN 0 0.054909f
C147 VIN 0 0.72895f
C148 sh_bsw3_1/ncell_bsw_sw_1/VBOOT 0 2.465944f
C149 CLKS 0 2.080142f
C150 sh_bsw3_0/cap_bsw_1/VPBT3 0 2.519834f
C151 sh_bsw3_0/cap_bsw_1/VPBT1 0 2.045305f
C152 sh_bsw3_0/cap_bsw_1/VPBT2 0 1.332593f
C153 sh_bsw3_0/ncell_bsw_dischrg_0/a_179_n1156# 0 0.084125f
C154 sh_bsw3_0/inv_bsw_0/VGND 0 1.846506f
C155 sh_bsw3_0/inv_bsw_0/OUT 0 0.977822f
C156 VCP 0 0.065191f
C157 VIP 0 0.741323f
C158 sh_bsw3_0/ncell_bsw_sw_1/VBOOT 0 2.465944f
.ends

