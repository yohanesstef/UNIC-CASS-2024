magic
tech sky130A
magscale 1 2
timestamp 1730722715
<< nwell >>
rect 611 -449 1297 145
<< nsubdiff >>
rect 647 75 749 109
rect 1159 75 1261 109
rect 647 17 681 75
rect 1227 17 1261 75
rect 647 -379 681 -325
rect 1227 -379 1261 -325
rect 647 -413 749 -379
rect 1159 -413 1261 -379
<< nsubdiffcont >>
rect 749 75 1159 109
rect 647 -325 681 17
rect 1227 -325 1261 17
rect 749 -413 1159 -379
<< poly >>
rect 807 -125 837 -109
rect 771 -135 837 -125
rect 771 -169 787 -135
rect 821 -169 837 -135
rect 771 -179 837 -169
rect 807 -199 837 -179
rect 895 -125 925 -109
rect 983 -125 1013 -109
rect 895 -135 1013 -125
rect 895 -169 925 -135
rect 983 -169 1013 -135
rect 895 -179 1013 -169
rect 895 -199 925 -179
rect 983 -199 1013 -179
rect 1071 -125 1101 -109
rect 1071 -135 1137 -125
rect 1071 -169 1087 -135
rect 1121 -169 1137 -135
rect 1071 -179 1137 -169
rect 1071 -199 1101 -179
<< polycont >>
rect 787 -169 821 -135
rect 925 -169 983 -135
rect 1087 -169 1121 -135
<< locali >>
rect 647 75 749 109
rect 1159 75 1261 109
rect 647 17 681 75
rect 761 21 795 75
rect 937 21 971 75
rect 1113 21 1147 75
rect 1227 17 1261 75
rect 761 -135 795 -87
rect 1113 -135 1147 -86
rect 761 -169 787 -135
rect 821 -169 837 -135
rect 909 -169 925 -135
rect 983 -169 999 -135
rect 1071 -169 1087 -135
rect 1121 -169 1147 -135
rect 761 -222 795 -169
rect 647 -379 681 -325
rect 761 -379 795 -327
rect 937 -379 971 -326
rect 1113 -379 1147 -169
rect 1227 -379 1261 -325
rect 647 -413 749 -379
rect 1159 -413 1261 -379
<< viali >>
rect 925 -169 983 -135
<< metal1 >>
rect 864 -1 892 17
rect 840 -7 892 -1
rect 840 -65 843 -59
rect 889 -65 892 -59
rect 1016 -1 1044 17
rect 1016 -7 1068 -1
rect 1016 -65 1068 -59
rect 925 -126 983 -123
rect 917 -135 991 -126
rect 917 -169 925 -135
rect 983 -169 991 -135
rect 917 -178 991 -169
rect 925 -181 983 -178
rect 840 -249 892 -243
rect 840 -307 892 -301
rect 1016 -249 1068 -243
rect 1016 -307 1068 -301
rect 861 -353 889 -320
rect 1019 -353 1047 -320
rect 861 -381 1047 -353
<< via1 >>
rect 840 -59 892 -7
rect 1016 -59 1068 -7
rect 840 -301 892 -249
rect 1016 -301 1068 -249
<< metal2 >>
rect 840 -7 892 -1
rect 840 -249 892 -59
rect 840 -307 892 -301
rect 1016 -7 1068 -1
rect 1016 -249 1068 -59
rect 1016 -307 1068 -301
use sky130_fd_pr__pfet_01v8_275TTJ  sky130_fd_pr__pfet_01v8_275TTJ_0
timestamp 1730448391
transform 1 0 910 0 1 -33
box -109 -112 109 112
use sky130_fd_pr__pfet_01v8_275TTJ  sky130_fd_pr__pfet_01v8_275TTJ_1
timestamp 1730448391
transform 1 0 998 0 1 -275
box -109 -112 109 112
use sky130_fd_pr__pfet_01v8_275TTJ  sky130_fd_pr__pfet_01v8_275TTJ_2
timestamp 1730448391
transform 1 0 910 0 1 -275
box -109 -112 109 112
use sky130_fd_pr__pfet_01v8_275TTJ  sky130_fd_pr__pfet_01v8_275TTJ_3
timestamp 1730448391
transform 1 0 822 0 1 -33
box -109 -112 109 112
use sky130_fd_pr__pfet_01v8_275TTJ  sky130_fd_pr__pfet_01v8_275TTJ_4
timestamp 1730448391
transform 1 0 1086 0 1 -33
box -109 -112 109 112
use sky130_fd_pr__pfet_01v8_275TTJ  sky130_fd_pr__pfet_01v8_275TTJ_6
timestamp 1730448391
transform 1 0 822 0 1 -275
box -109 -112 109 112
use sky130_fd_pr__pfet_01v8_275TTJ  sky130_fd_pr__pfet_01v8_275TTJ_7
timestamp 1730448391
transform 1 0 998 0 1 -33
box -109 -112 109 112
use sky130_fd_pr__pfet_01v8_275TTJ  sky130_fd_pr__pfet_01v8_275TTJ_8
timestamp 1730448391
transform 1 0 1086 0 1 -275
box -109 -112 109 112
<< labels >>
flabel viali 954 -152 954 -152 0 FreeSans 80 0 0 0 SWITCHING
port 2 nsew
flabel metal2 s 866 -275 866 -275 0 FreeSans 80 0 0 0 VBOOT
port 3 nsew
flabel locali s 954 92 954 92 0 FreeSans 320 0 0 0 VPBT3
port 1 nsew
<< end >>
