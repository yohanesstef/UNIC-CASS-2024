magic
tech sky130A
magscale 1 2
timestamp 1730800698
<< nwell >>
rect 1301 216 1439 262
<< pwell >>
rect 2689 2110 2741 2116
rect 2683 2058 2747 2110
rect 2683 990 2747 1042
rect 3795 809 3991 875
<< locali >>
rect 1561 2225 1757 2291
rect 3795 809 3991 875
rect 3431 350 3625 530
rect 3431 282 3437 350
rect 3619 282 3625 350
rect 3431 276 3625 282
<< viali >>
rect 4205 2768 4239 2866
rect 1313 234 1347 332
rect 3437 282 3619 350
<< metal1 >>
rect 1277 3102 1678 3258
rect 1730 3102 3906 3258
rect 3958 3102 4275 3258
rect 4129 2866 4251 2884
rect 4129 2838 4205 2866
rect 4193 2768 4205 2838
rect 4239 2768 4251 2866
rect 4193 2761 4251 2768
rect 1672 2232 1678 2284
rect 2683 2058 2689 2110
rect 2741 2058 2747 2110
rect 2683 990 2689 1042
rect 2741 990 2747 1042
rect 3795 861 3875 875
rect 3795 809 3817 861
rect 3869 809 3875 861
rect 3431 350 3625 362
rect 1301 332 1359 339
rect 1301 234 1313 332
rect 1347 262 1359 332
rect 3431 282 3437 350
rect 3619 282 3625 350
rect 3431 270 3625 282
rect 1347 234 1439 262
rect 1301 216 1439 234
rect 1277 -158 3431 -2
rect 3625 -158 4275 -2
<< via1 >>
rect 1678 3102 1730 3258
rect 3906 3102 3958 3258
rect 1678 2232 1730 2284
rect 2689 2058 2741 2110
rect 2689 990 2741 1042
rect 3817 809 3869 861
rect 3437 282 3619 350
rect 3431 -158 3625 -2
<< metal2 >>
rect 1678 3258 1730 3264
rect 1678 2284 1730 3102
rect 3906 3258 3958 3264
rect 3906 2702 3958 3102
rect 1678 1866 1730 2232
rect 1594 1814 1730 1866
rect 2689 2110 2741 2116
rect 1594 1425 1646 1814
rect 2689 1042 2741 2058
rect 2811 1997 2871 2006
rect 2811 1162 2871 1937
rect 3906 1283 3958 1669
rect 3817 1231 3958 1283
rect 2804 1106 2813 1162
rect 2869 1106 2878 1162
rect 2811 1104 2871 1106
rect 2689 984 2741 990
rect 3817 861 3869 1231
rect 3817 803 3869 809
rect 3431 350 3625 357
rect 3431 282 3437 350
rect 3619 282 3625 350
rect 3431 -2 3625 282
rect 3431 -164 3625 -158
<< via2 >>
rect 2811 1937 2871 1997
rect 2813 1106 2869 1162
<< metal3 >>
rect 2806 1997 2876 2002
rect 2806 1937 2811 1997
rect 2871 1937 4412 1997
rect 2806 1932 2876 1937
rect 2808 1164 2874 1167
rect 1177 1162 2874 1164
rect 1177 1106 2813 1162
rect 2869 1106 2874 1162
rect 1177 1104 2874 1106
rect 2808 1101 2874 1104
use sh_bsw3  sh_bsw3_0
timestamp 1730800306
transform -1 0 4275 0 -1 2708
box -1300 -376 2998 1784
use sh_bsw3  sh_bsw3_1
timestamp 1730800306
transform 1 0 1277 0 1 392
box -1300 -376 2998 1784
<< labels >>
flabel metal1 s 1277 3182 1277 3182 3 FreeSans 480 0 0 0 VDDA
port 1 e
flabel metal1 s 1201 154 1201 154 3 FreeSans 480 0 0 0 CLKS
port 2 e
flabel metal1 s 1201 49 1201 49 3 FreeSans 480 0 0 0 CLKSB
port 3 e
flabel metal2 s 2655 2808 2655 2808 3 FreeSans 480 0 0 0 VIP
port 4 e
flabel metal2 s 2657 291 2657 291 3 FreeSans 480 0 0 0 VIN
port 5 e
flabel metal1 s 1277 -95 1277 -95 3 FreeSans 480 0 0 0 VSSA
port 6 e
flabel metal2 s 2776 2934 2776 2934 0 FreeSans 480 0 0 0 VCP
port 7 nsew
flabel metal2 s 2776 164 2776 164 0 FreeSans 480 0 0 0 VCN
port 8 nsew
<< end >>
