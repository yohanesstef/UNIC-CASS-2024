magic
tech sky130A
magscale 1 2
timestamp 1730612622
<< pwell >>
rect -567 -3799 943 -2748
<< ndiff >>
rect -186 -3172 -134 -3120
rect 510 -3172 562 -3120
rect 598 -3172 650 -3120
rect -186 -3427 -134 -3375
rect 510 -3427 562 -3375
<< psubdiff >>
rect -531 -2818 -417 -2784
rect 793 -2818 907 -2784
rect -531 -2870 -497 -2818
rect 873 -2870 907 -2818
rect -531 -3729 -497 -3604
rect 873 -3729 907 -3604
rect -531 -3763 -417 -3729
rect 793 -3763 907 -3729
<< psubdiffcont >>
rect -417 -2818 793 -2784
rect -531 -3604 -497 -2870
rect 873 -3604 907 -2870
rect -417 -3763 793 -3729
<< poly >>
rect 335 -3024 401 -3008
rect 335 -3058 351 -3024
rect 385 -3058 401 -3024
rect 335 -3074 401 -3058
rect 529 -3024 595 -3009
rect 529 -3058 545 -3024
rect 579 -3058 595 -3024
rect 529 -3075 595 -3058
rect 653 -3024 719 -3008
rect 653 -3058 669 -3024
rect 703 -3058 719 -3024
rect 653 -3074 719 -3058
rect -343 -3234 -277 -3218
rect -343 -3268 -327 -3234
rect -293 -3268 -277 -3234
rect -343 -3284 -277 -3268
rect -219 -3234 -153 -3218
rect -219 -3268 -203 -3234
rect -169 -3268 -153 -3234
rect -219 -3284 -153 -3268
rect -19 -3234 47 -3218
rect -19 -3268 -3 -3234
rect 31 -3268 47 -3234
rect -19 -3284 47 -3268
rect 99 -3234 159 -3222
rect 99 -3268 112 -3234
rect 146 -3268 159 -3234
rect 99 -3326 159 -3268
rect 217 -3280 277 -3222
rect 217 -3314 230 -3280
rect 264 -3314 277 -3280
rect 217 -3326 277 -3314
rect 329 -3280 395 -3264
rect 329 -3314 345 -3280
rect 379 -3314 395 -3280
rect 329 -3330 395 -3314
rect 529 -3280 595 -3264
rect 529 -3314 545 -3280
rect 579 -3314 595 -3280
rect 529 -3330 595 -3314
rect 653 -3280 719 -3264
rect 653 -3314 669 -3280
rect 703 -3314 719 -3280
rect 653 -3330 719 -3314
rect -343 -3490 -277 -3474
rect -343 -3524 -327 -3490
rect -293 -3524 -277 -3490
rect -343 -3540 -277 -3524
rect -219 -3490 -153 -3474
rect -219 -3524 -203 -3490
rect -169 -3524 -153 -3490
rect -219 -3540 -153 -3524
rect -25 -3490 41 -3474
rect -25 -3524 -9 -3490
rect 25 -3524 41 -3490
rect -25 -3540 41 -3524
<< polycont >>
rect 351 -3058 385 -3024
rect 545 -3058 579 -3024
rect 669 -3058 703 -3024
rect -327 -3268 -293 -3234
rect -203 -3268 -169 -3234
rect -3 -3268 31 -3234
rect 112 -3268 146 -3234
rect 230 -3314 264 -3280
rect 345 -3314 379 -3280
rect 545 -3314 579 -3280
rect 669 -3314 703 -3280
rect -327 -3524 -293 -3490
rect -203 -3524 -169 -3490
rect -9 -3524 25 -3490
<< locali >>
rect -531 -2818 -417 -2784
rect 793 -2818 907 -2784
rect -531 -2870 -497 -2818
rect 873 -2870 907 -2818
rect 335 -3058 351 -3024
rect 385 -3058 401 -3024
rect 529 -3058 545 -3024
rect 579 -3058 595 -3024
rect 653 -3058 669 -3024
rect 703 -3058 719 -3024
rect -343 -3268 -327 -3234
rect -293 -3268 -277 -3234
rect -219 -3268 -203 -3234
rect -169 -3268 -153 -3234
rect -19 -3268 -3 -3234
rect 31 -3268 47 -3234
rect 96 -3268 112 -3234
rect 146 -3268 162 -3234
rect 214 -3314 230 -3280
rect 264 -3314 280 -3280
rect 329 -3314 345 -3280
rect 379 -3314 395 -3280
rect 529 -3314 545 -3280
rect 579 -3314 595 -3280
rect 653 -3314 669 -3280
rect 703 -3314 719 -3280
rect -343 -3524 -327 -3490
rect -293 -3524 -277 -3490
rect -219 -3524 -203 -3490
rect -169 -3524 -153 -3490
rect -25 -3524 -9 -3490
rect 25 -3524 41 -3490
rect -531 -3729 -497 -3604
rect 873 -3729 907 -3604
rect -531 -3763 -417 -3729
rect 793 -3763 907 -3729
<< viali >>
rect 351 -3058 385 -3024
rect 545 -3058 579 -3024
rect 669 -3058 703 -3024
rect 866 -3058 873 -3024
rect 873 -3058 900 -3024
rect -327 -3268 -293 -3234
rect -203 -3268 -169 -3234
rect -3 -3268 31 -3234
rect 112 -3268 146 -3234
rect 230 -3314 264 -3280
rect 345 -3314 379 -3280
rect 545 -3314 579 -3280
rect 669 -3314 703 -3280
rect -525 -3524 -497 -3490
rect -497 -3524 -491 -3490
rect -327 -3524 -293 -3490
rect -203 -3524 -169 -3490
rect -9 -3524 25 -3490
<< metal1 >>
rect -497 -2877 793 -2870
rect -445 -2916 741 -2877
rect -497 -2935 -445 -2929
rect 741 -2935 793 -2929
rect -417 -2950 585 -2944
rect -365 -2990 585 -2950
rect -417 -3008 -365 -3002
rect 345 -3022 391 -3018
rect 47 -3024 447 -3022
rect 539 -3024 585 -2990
rect 873 -3018 907 -3012
rect 619 -3024 907 -3018
rect 47 -3058 351 -3024
rect 385 -3058 447 -3024
rect 533 -3058 545 -3024
rect 579 -3058 591 -3024
rect 619 -3058 669 -3024
rect 703 -3058 866 -3024
rect 900 -3058 907 -3024
rect 47 -3064 447 -3058
rect 539 -3064 585 -3058
rect 619 -3064 907 -3058
rect 47 -3068 329 -3064
rect 47 -3096 93 -3068
rect 283 -3096 329 -3068
rect -183 -3114 -25 -3096
rect 401 -3100 447 -3064
rect 619 -3096 647 -3064
rect 689 -3096 735 -3064
rect 873 -3070 907 -3064
rect -186 -3120 -25 -3114
rect -134 -3172 -25 -3120
rect -186 -3178 -25 -3172
rect 44 -3120 96 -3114
rect 44 -3178 96 -3172
rect 162 -3120 214 -3114
rect 162 -3178 214 -3172
rect 280 -3120 332 -3114
rect 280 -3178 332 -3172
rect 510 -3120 562 -3114
rect 510 -3178 562 -3172
rect -497 -3207 -445 -3201
rect -359 -3228 -313 -3196
rect -271 -3228 -243 -3184
rect -183 -3196 -25 -3178
rect -359 -3234 -243 -3228
rect -209 -3234 -163 -3228
rect -9 -3234 37 -3228
rect 106 -3234 152 -3228
rect -445 -3259 -327 -3234
rect -497 -3268 -327 -3259
rect -293 -3268 -243 -3234
rect -215 -3268 -203 -3234
rect -169 -3268 -3 -3234
rect 31 -3268 112 -3234
rect 146 -3268 270 -3234
rect -359 -3274 -243 -3268
rect -209 -3274 -163 -3268
rect -9 -3274 37 -3268
rect 106 -3280 270 -3268
rect 741 -3262 793 -3256
rect 339 -3280 385 -3274
rect 539 -3280 585 -3274
rect 619 -3280 741 -3274
rect 106 -3314 230 -3280
rect 264 -3314 345 -3280
rect 379 -3314 545 -3280
rect 579 -3314 591 -3280
rect 619 -3314 669 -3280
rect 703 -3314 741 -3280
rect 224 -3320 270 -3314
rect 339 -3320 385 -3314
rect 539 -3320 585 -3314
rect 619 -3320 793 -3314
rect 401 -3369 559 -3352
rect 619 -3364 647 -3320
rect 689 -3352 735 -3320
rect -186 -3375 -134 -3369
rect -186 -3433 -134 -3427
rect 44 -3375 96 -3369
rect 44 -3433 96 -3427
rect 162 -3375 214 -3369
rect 162 -3433 214 -3427
rect 280 -3375 332 -3369
rect 280 -3433 332 -3427
rect 401 -3375 562 -3369
rect 401 -3427 510 -3375
rect 401 -3433 562 -3427
rect -531 -3484 -497 -3478
rect -359 -3484 -313 -3440
rect -271 -3484 -243 -3440
rect 401 -3452 559 -3433
rect -71 -3480 -25 -3452
rect 47 -3480 93 -3452
rect 283 -3480 329 -3452
rect -531 -3490 -243 -3484
rect -531 -3524 -525 -3490
rect -491 -3524 -327 -3490
rect -293 -3524 -243 -3490
rect -531 -3530 -243 -3524
rect -215 -3490 -157 -3480
rect -215 -3524 -203 -3490
rect -169 -3524 -157 -3490
rect -215 -3530 -157 -3524
rect -71 -3490 329 -3480
rect -71 -3524 -9 -3490
rect 25 -3524 329 -3490
rect -71 -3526 329 -3524
rect -15 -3530 31 -3526
rect -531 -3536 -497 -3530
rect -209 -3558 -163 -3530
rect 510 -3546 562 -3540
rect -423 -3610 -417 -3558
rect -365 -3604 -163 -3558
rect -365 -3610 -359 -3604
rect -83 -3610 -77 -3558
rect -25 -3598 510 -3558
rect -25 -3604 562 -3598
rect -25 -3610 -19 -3604
<< via1 >>
rect -497 -2929 -445 -2877
rect 741 -2929 793 -2877
rect -417 -3002 -365 -2950
rect -186 -3172 -134 -3120
rect 44 -3172 96 -3120
rect 162 -3172 214 -3120
rect 280 -3172 332 -3120
rect 510 -3172 562 -3120
rect -497 -3259 -445 -3207
rect 741 -3314 793 -3262
rect -186 -3427 -134 -3375
rect 44 -3427 96 -3375
rect 162 -3427 214 -3375
rect 280 -3427 332 -3375
rect 510 -3427 562 -3375
rect -417 -3610 -365 -3558
rect -77 -3610 -25 -3558
rect 510 -3598 562 -3546
<< metal2 >>
rect -497 -2877 -445 -2870
rect -497 -3207 -445 -2929
rect 741 -2877 793 -2870
rect -497 -3268 -445 -3259
rect -417 -2950 -365 -2944
rect -417 -3558 -365 -3002
rect -186 -3120 -134 -3114
rect -186 -3375 -134 -3172
rect -186 -3558 -134 -3427
rect 44 -3120 96 -3114
rect 44 -3375 96 -3172
rect 44 -3433 96 -3427
rect 162 -3120 214 -3114
rect 162 -3375 214 -3172
rect 162 -3433 214 -3427
rect 280 -3120 332 -3114
rect 280 -3375 332 -3172
rect 280 -3433 332 -3427
rect 510 -3120 562 -3114
rect 510 -3375 562 -3172
rect 741 -3262 793 -2929
rect 741 -3320 793 -3314
rect 510 -3546 562 -3427
rect -186 -3604 -77 -3558
rect -83 -3610 -77 -3604
rect -25 -3610 -19 -3558
rect 510 -3604 562 -3598
rect -417 -3616 -365 -3610
use sky130_fd_pr__nfet_01v8_6J3TAM  sky130_fd_pr__nfet_01v8_6J3TAM_0
timestamp 1730478237
transform 1 0 -204 0 1 -3146
box -73 -76 73 76
use sky130_fd_pr__nfet_01v8_6J3TAM  sky130_fd_pr__nfet_01v8_6J3TAM_1
timestamp 1730478237
transform 1 0 580 0 1 -3402
box -73 -76 73 76
use sky130_fd_pr__nfet_01v8_6J3TAM  sky130_fd_pr__nfet_01v8_6J3TAM_2
timestamp 1730478237
transform 1 0 -204 0 1 -3402
box -73 -76 73 76
use sky130_fd_pr__nfet_01v8_6J3TAM  sky130_fd_pr__nfet_01v8_6J3TAM_3
timestamp 1730478237
transform 1 0 580 0 1 -3146
box -73 -76 73 76
use sky130_fd_pr__nfet_01v8_6J3TAM  sky130_fd_pr__nfet_01v8_6J3TAM_4
timestamp 1730478237
transform 1 0 668 0 1 -3146
box -73 -76 73 76
use sky130_fd_pr__nfet_01v8_6J3TAM  sky130_fd_pr__nfet_01v8_6J3TAM_5
timestamp 1730478237
transform 1 0 -292 0 1 -3402
box -73 -76 73 76
use sky130_fd_pr__nfet_01v8_6J3TAM  sky130_fd_pr__nfet_01v8_6J3TAM_6
timestamp 1730478237
transform 1 0 668 0 1 -3402
box -73 -76 73 76
use sky130_fd_pr__nfet_01v8_6J3TAM  sky130_fd_pr__nfet_01v8_6J3TAM_10
timestamp 1730478237
transform 1 0 -292 0 1 -3146
box -73 -76 73 76
use sky130_fd_pr__nfet_01v8_QS6TK8  sky130_fd_pr__nfet_01v8_QS6TK8_0
timestamp 1730569521
transform 1 0 11 0 1 -3146
box -88 -76 88 76
use sky130_fd_pr__nfet_01v8_QS6TK8  sky130_fd_pr__nfet_01v8_QS6TK8_1
timestamp 1730569521
transform 1 0 129 0 1 -3146
box -88 -76 88 76
use sky130_fd_pr__nfet_01v8_QS6TK8  sky130_fd_pr__nfet_01v8_QS6TK8_2
timestamp 1730569521
transform 1 0 247 0 1 -3146
box -88 -76 88 76
use sky130_fd_pr__nfet_01v8_QS6TK8  sky130_fd_pr__nfet_01v8_QS6TK8_3
timestamp 1730569521
transform 1 0 365 0 1 -3402
box -88 -76 88 76
use sky130_fd_pr__nfet_01v8_QS6TK8  sky130_fd_pr__nfet_01v8_QS6TK8_4
timestamp 1730569521
transform 1 0 365 0 1 -3146
box -88 -76 88 76
use sky130_fd_pr__nfet_01v8_QS6TK8  sky130_fd_pr__nfet_01v8_QS6TK8_5
timestamp 1730569521
transform 1 0 11 0 1 -3402
box -88 -76 88 76
use sky130_fd_pr__nfet_01v8_QS6TK8  sky130_fd_pr__nfet_01v8_QS6TK8_6
timestamp 1730569521
transform 1 0 129 0 1 -3402
box -88 -76 88 76
use sky130_fd_pr__nfet_01v8_QS6TK8  sky130_fd_pr__nfet_01v8_QS6TK8_7
timestamp 1730569521
transform 1 0 247 0 1 -3402
box -88 -76 88 76
<< labels >>
flabel metal1 s -73 -3251 -73 -3251 0 FreeSans 240 0 0 0 VBOOT
port 2 nsew
flabel metal1 s 117 -2966 117 -2966 0 FreeSans 240 0 0 0 VNBT1
port 3 nsew
flabel metal1 s 216 -3582 216 -3582 0 FreeSans 240 0 0 0 VNBT3
port 4 nsew
flabel metal1 s 112 -2891 112 -2891 0 FreeSans 240 0 0 0 SWITCHING
port 5 nsew
flabel locali s 158 -2801 158 -2801 0 FreeSans 240 0 0 0 VSSA
port 6 nsew
flabel metal2 s 188 -3212 188 -3212 0 FreeSans 240 0 0 0 VO
port 7 nsew
flabel metal1 s 190 -3506 190 -3506 0 FreeSans 240 0 0 0 VI
port 1 nsew
<< end >>
